// testbench_ls.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module testbench_ls (
		output wire         clk_200_out_clk_clk,                                     //                              clk_200_out_clk.clk
		input  wire         clk_50_clk,                                              //                                       clk_50.clk
		output wire [3:0]   ctrl_sig_export,                                         //                                     ctrl_sig.export
		output wire         ddr2_ram_status_local_init_done,                         //                              ddr2_ram_status.local_init_done
		output wire         ddr2_ram_status_local_cal_success,                       //                                             .local_cal_success
		output wire         ddr2_ram_status_local_cal_fail,                          //                                             .local_cal_fail
		output wire [255:0] dma_fifo_subsystem_2_fifo_stream_conduit_end_fifo_data,  // dma_fifo_subsystem_2_fifo_stream_conduit_end.fifo_data
		output wire         dma_fifo_subsystem_2_fifo_stream_conduit_end_fifo_write, //                                             .fifo_write
		output wire         dma_fifo_subsystem_2_fifo_stream_conduit_end_fifo_send,  //                                             .fifo_send
		output wire [255:0] dma_fifo_subsystem_3_fifo_stream_conduit_end_fifo_data,  // dma_fifo_subsystem_3_fifo_stream_conduit_end.fifo_data
		output wire         dma_fifo_subsystem_3_fifo_stream_conduit_end_fifo_write, //                                             .fifo_write
		output wire         dma_fifo_subsystem_3_fifo_stream_conduit_end_fifo_send,  //                                             .fifo_send
		output wire [255:0] dma_fifo_subsystem_4_fifo_stream_conduit_end_fifo_data,  // dma_fifo_subsystem_4_fifo_stream_conduit_end.fifo_data
		output wire         dma_fifo_subsystem_4_fifo_stream_conduit_end_fifo_write, //                                             .fifo_write
		output wire         dma_fifo_subsystem_4_fifo_stream_conduit_end_fifo_send,  //                                             .fifo_send
		output wire [255:0] fifo_stream_fifo_data,                                   //                                  fifo_stream.fifo_data
		output wire         fifo_stream_fifo_write,                                  //                                             .fifo_write
		output wire         fifo_stream_fifo_send,                                   //                                             .fifo_send
		output wire [255:0] fifo_stream_1_fifo_data,                                 //                                fifo_stream_1.fifo_data
		output wire         fifo_stream_1_fifo_write,                                //                                             .fifo_write
		output wire         fifo_stream_1_fifo_send,                                 //                                             .fifo_send
		input  wire [63:0]  from_fifo_fifo_data,                                     //                                    from_fifo.fifo_data
		output wire         from_fifo_fifo_read,                                     //                                             .fifo_read
		input  wire         from_fifo_fifo_empty,                                    //                                             .fifo_empty
		input  wire         from_fifo_fifo_full,                                     //                                             .fifo_full
		input  wire [15:0]  input_io_0_external_connection_export,                   //               input_io_0_external_connection.export
		input  wire [15:0]  input_io_1_external_connection_export,                   //               input_io_1_external_connection.export
		input  wire [15:0]  input_io_2_external_connection_export,                   //               input_io_2_external_connection.export
		input  wire [15:0]  input_io_3_external_connection_export,                   //               input_io_3_external_connection.export
		input  wire [15:0]  input_io_4_external_connection_export,                   //               input_io_4_external_connection.export
		input  wire [7:0]   input_io_5_external_connection_export,                   //               input_io_5_external_connection.export
		input  wire [15:0]  input_io_external_connection_export,                     //                 input_io_external_connection.export
		output wire [13:0]  memory_mem_a,                                            //                                       memory.mem_a
		output wire [2:0]   memory_mem_ba,                                           //                                             .mem_ba
		output wire [1:0]   memory_mem_ck,                                           //                                             .mem_ck
		output wire [1:0]   memory_mem_ck_n,                                         //                                             .mem_ck_n
		output wire [0:0]   memory_mem_cke,                                          //                                             .mem_cke
		output wire [0:0]   memory_mem_cs_n,                                         //                                             .mem_cs_n
		output wire [7:0]   memory_mem_dm,                                           //                                             .mem_dm
		output wire [0:0]   memory_mem_ras_n,                                        //                                             .mem_ras_n
		output wire [0:0]   memory_mem_cas_n,                                        //                                             .mem_cas_n
		output wire [0:0]   memory_mem_we_n,                                         //                                             .mem_we_n
		inout  wire [63:0]  memory_mem_dq,                                           //                                             .mem_dq
		inout  wire [7:0]   memory_mem_dqs,                                          //                                             .mem_dqs
		inout  wire [7:0]   memory_mem_dqs_n,                                        //                                             .mem_dqs_n
		output wire [0:0]   memory_mem_odt,                                          //                                             .mem_odt
		output wire [13:0]  memory_1_mem_a,                                          //                                     memory_1.mem_a
		output wire [2:0]   memory_1_mem_ba,                                         //                                             .mem_ba
		output wire [1:0]   memory_1_mem_ck,                                         //                                             .mem_ck
		output wire [1:0]   memory_1_mem_ck_n,                                       //                                             .mem_ck_n
		output wire [0:0]   memory_1_mem_cke,                                        //                                             .mem_cke
		output wire [0:0]   memory_1_mem_cs_n,                                       //                                             .mem_cs_n
		output wire [7:0]   memory_1_mem_dm,                                         //                                             .mem_dm
		output wire [0:0]   memory_1_mem_ras_n,                                      //                                             .mem_ras_n
		output wire [0:0]   memory_1_mem_cas_n,                                      //                                             .mem_cas_n
		output wire [0:0]   memory_1_mem_we_n,                                       //                                             .mem_we_n
		inout  wire [63:0]  memory_1_mem_dq,                                         //                                             .mem_dq
		inout  wire [7:0]   memory_1_mem_dqs,                                        //                                             .mem_dqs
		inout  wire [7:0]   memory_1_mem_dqs_n,                                      //                                             .mem_dqs_n
		output wire [0:0]   memory_1_mem_odt,                                        //                                             .mem_odt
		input  wire         oct_rdn,                                                 //                                          oct.rdn
		input  wire         oct_rup,                                                 //                                             .rup
		input  wire         oct_1_rdn,                                               //                                        oct_1.rdn
		input  wire         oct_1_rup,                                               //                                             .rup
		input  wire [7:0]   pilot_sig_external_connection_export,                    //                pilot_sig_external_connection.export
		input  wire         reset_reset_n                                            //                                        reset.reset_n
	);

	wire          from_eth_to_ddr_eth_dma_mm_write_waitrequest;                            // mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_mm_write_waitrequest -> from_ETH_to_DDR:ETH_DMA_mm_write_waitrequest
	wire   [30:0] from_eth_to_ddr_eth_dma_mm_write_address;                                // from_ETH_to_DDR:ETH_DMA_mm_write_address -> mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_mm_write_address
	wire   [31:0] from_eth_to_ddr_eth_dma_mm_write_byteenable;                             // from_ETH_to_DDR:ETH_DMA_mm_write_byteenable -> mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_mm_write_byteenable
	wire          from_eth_to_ddr_eth_dma_mm_write_write;                                  // from_ETH_to_DDR:ETH_DMA_mm_write_write -> mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_mm_write_write
	wire  [255:0] from_eth_to_ddr_eth_dma_mm_write_writedata;                              // from_ETH_to_DDR:ETH_DMA_mm_write_writedata -> mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_mm_write_writedata
	wire   [31:0] nios_cpu_data_master_readdata;                                           // mm_interconnect_0:nios_cpu_data_master_readdata -> nios_cpu:d_readdata
	wire          nios_cpu_data_master_waitrequest;                                        // mm_interconnect_0:nios_cpu_data_master_waitrequest -> nios_cpu:d_waitrequest
	wire          nios_cpu_data_master_debugaccess;                                        // nios_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_cpu_data_master_debugaccess
	wire   [31:0] nios_cpu_data_master_address;                                            // nios_cpu:d_address -> mm_interconnect_0:nios_cpu_data_master_address
	wire    [3:0] nios_cpu_data_master_byteenable;                                         // nios_cpu:d_byteenable -> mm_interconnect_0:nios_cpu_data_master_byteenable
	wire          nios_cpu_data_master_read;                                               // nios_cpu:d_read -> mm_interconnect_0:nios_cpu_data_master_read
	wire          nios_cpu_data_master_readdatavalid;                                      // mm_interconnect_0:nios_cpu_data_master_readdatavalid -> nios_cpu:d_readdatavalid
	wire          nios_cpu_data_master_write;                                              // nios_cpu:d_write -> mm_interconnect_0:nios_cpu_data_master_write
	wire   [31:0] nios_cpu_data_master_writedata;                                          // nios_cpu:d_writedata -> mm_interconnect_0:nios_cpu_data_master_writedata
	wire  [255:0] dma_fifo_susbystem_dma_mm_read_readdata;                                 // mm_interconnect_0:dma_fifo_susbystem_dma_mm_read_readdata -> dma_fifo_susbystem:dma_mm_read_readdata
	wire          dma_fifo_susbystem_dma_mm_read_waitrequest;                              // mm_interconnect_0:dma_fifo_susbystem_dma_mm_read_waitrequest -> dma_fifo_susbystem:dma_mm_read_waitrequest
	wire   [29:0] dma_fifo_susbystem_dma_mm_read_address;                                  // dma_fifo_susbystem:dma_mm_read_address -> mm_interconnect_0:dma_fifo_susbystem_dma_mm_read_address
	wire          dma_fifo_susbystem_dma_mm_read_read;                                     // dma_fifo_susbystem:dma_mm_read_read -> mm_interconnect_0:dma_fifo_susbystem_dma_mm_read_read
	wire   [31:0] dma_fifo_susbystem_dma_mm_read_byteenable;                               // dma_fifo_susbystem:dma_mm_read_byteenable -> mm_interconnect_0:dma_fifo_susbystem_dma_mm_read_byteenable
	wire          dma_fifo_susbystem_dma_mm_read_readdatavalid;                            // mm_interconnect_0:dma_fifo_susbystem_dma_mm_read_readdatavalid -> dma_fifo_susbystem:dma_mm_read_readdatavalid
	wire   [10:0] dma_fifo_susbystem_dma_mm_read_burstcount;                               // dma_fifo_susbystem:dma_mm_read_burstcount -> mm_interconnect_0:dma_fifo_susbystem_dma_mm_read_burstcount
	wire  [255:0] dma_fifo_subsystem_1_dma_mm_read_readdata;                               // mm_interconnect_0:dma_fifo_subsystem_1_dma_mm_read_readdata -> dma_fifo_subsystem_1:dma_mm_read_readdata
	wire          dma_fifo_subsystem_1_dma_mm_read_waitrequest;                            // mm_interconnect_0:dma_fifo_subsystem_1_dma_mm_read_waitrequest -> dma_fifo_subsystem_1:dma_mm_read_waitrequest
	wire   [29:0] dma_fifo_subsystem_1_dma_mm_read_address;                                // dma_fifo_subsystem_1:dma_mm_read_address -> mm_interconnect_0:dma_fifo_subsystem_1_dma_mm_read_address
	wire          dma_fifo_subsystem_1_dma_mm_read_read;                                   // dma_fifo_subsystem_1:dma_mm_read_read -> mm_interconnect_0:dma_fifo_subsystem_1_dma_mm_read_read
	wire   [31:0] dma_fifo_subsystem_1_dma_mm_read_byteenable;                             // dma_fifo_subsystem_1:dma_mm_read_byteenable -> mm_interconnect_0:dma_fifo_subsystem_1_dma_mm_read_byteenable
	wire          dma_fifo_subsystem_1_dma_mm_read_readdatavalid;                          // mm_interconnect_0:dma_fifo_subsystem_1_dma_mm_read_readdatavalid -> dma_fifo_subsystem_1:dma_mm_read_readdatavalid
	wire   [10:0] dma_fifo_subsystem_1_dma_mm_read_burstcount;                             // dma_fifo_subsystem_1:dma_mm_read_burstcount -> mm_interconnect_0:dma_fifo_subsystem_1_dma_mm_read_burstcount
	wire  [255:0] dma_fifo_subsystem_2_dma_mm_read_readdata;                               // mm_interconnect_0:dma_fifo_subsystem_2_dma_mm_read_readdata -> dma_fifo_subsystem_2:dma_mm_read_readdata
	wire          dma_fifo_subsystem_2_dma_mm_read_waitrequest;                            // mm_interconnect_0:dma_fifo_subsystem_2_dma_mm_read_waitrequest -> dma_fifo_subsystem_2:dma_mm_read_waitrequest
	wire   [29:0] dma_fifo_subsystem_2_dma_mm_read_address;                                // dma_fifo_subsystem_2:dma_mm_read_address -> mm_interconnect_0:dma_fifo_subsystem_2_dma_mm_read_address
	wire          dma_fifo_subsystem_2_dma_mm_read_read;                                   // dma_fifo_subsystem_2:dma_mm_read_read -> mm_interconnect_0:dma_fifo_subsystem_2_dma_mm_read_read
	wire   [31:0] dma_fifo_subsystem_2_dma_mm_read_byteenable;                             // dma_fifo_subsystem_2:dma_mm_read_byteenable -> mm_interconnect_0:dma_fifo_subsystem_2_dma_mm_read_byteenable
	wire          dma_fifo_subsystem_2_dma_mm_read_readdatavalid;                          // mm_interconnect_0:dma_fifo_subsystem_2_dma_mm_read_readdatavalid -> dma_fifo_subsystem_2:dma_mm_read_readdatavalid
	wire   [10:0] dma_fifo_subsystem_2_dma_mm_read_burstcount;                             // dma_fifo_subsystem_2:dma_mm_read_burstcount -> mm_interconnect_0:dma_fifo_subsystem_2_dma_mm_read_burstcount
	wire   [31:0] nios_cpu_instruction_master_readdata;                                    // mm_interconnect_0:nios_cpu_instruction_master_readdata -> nios_cpu:i_readdata
	wire          nios_cpu_instruction_master_waitrequest;                                 // mm_interconnect_0:nios_cpu_instruction_master_waitrequest -> nios_cpu:i_waitrequest
	wire   [31:0] nios_cpu_instruction_master_address;                                     // nios_cpu:i_address -> mm_interconnect_0:nios_cpu_instruction_master_address
	wire          nios_cpu_instruction_master_read;                                        // nios_cpu:i_read -> mm_interconnect_0:nios_cpu_instruction_master_read
	wire          nios_cpu_instruction_master_readdatavalid;                               // mm_interconnect_0:nios_cpu_instruction_master_readdatavalid -> nios_cpu:i_readdatavalid
	wire  [255:0] dma_fifo_subsystem_4_dma_mm_read_readdata;                               // mm_interconnect_0:dma_fifo_subsystem_4_dma_mm_read_readdata -> dma_fifo_subsystem_4:dma_mm_read_readdata
	wire          dma_fifo_subsystem_4_dma_mm_read_waitrequest;                            // mm_interconnect_0:dma_fifo_subsystem_4_dma_mm_read_waitrequest -> dma_fifo_subsystem_4:dma_mm_read_waitrequest
	wire   [30:0] dma_fifo_subsystem_4_dma_mm_read_address;                                // dma_fifo_subsystem_4:dma_mm_read_address -> mm_interconnect_0:dma_fifo_subsystem_4_dma_mm_read_address
	wire          dma_fifo_subsystem_4_dma_mm_read_read;                                   // dma_fifo_subsystem_4:dma_mm_read_read -> mm_interconnect_0:dma_fifo_subsystem_4_dma_mm_read_read
	wire   [31:0] dma_fifo_subsystem_4_dma_mm_read_byteenable;                             // dma_fifo_subsystem_4:dma_mm_read_byteenable -> mm_interconnect_0:dma_fifo_subsystem_4_dma_mm_read_byteenable
	wire          dma_fifo_subsystem_4_dma_mm_read_readdatavalid;                          // mm_interconnect_0:dma_fifo_subsystem_4_dma_mm_read_readdatavalid -> dma_fifo_subsystem_4:dma_mm_read_readdatavalid
	wire   [10:0] dma_fifo_subsystem_4_dma_mm_read_burstcount;                             // dma_fifo_subsystem_4:dma_mm_read_burstcount -> mm_interconnect_0:dma_fifo_subsystem_4_dma_mm_read_burstcount
	wire  [255:0] dma_fifo_subsystem_3_dma_mm_read_readdata;                               // mm_interconnect_0:dma_fifo_subsystem_3_dma_mm_read_readdata -> dma_fifo_subsystem_3:dma_mm_read_readdata
	wire          dma_fifo_subsystem_3_dma_mm_read_waitrequest;                            // mm_interconnect_0:dma_fifo_subsystem_3_dma_mm_read_waitrequest -> dma_fifo_subsystem_3:dma_mm_read_waitrequest
	wire   [30:0] dma_fifo_subsystem_3_dma_mm_read_address;                                // dma_fifo_subsystem_3:dma_mm_read_address -> mm_interconnect_0:dma_fifo_subsystem_3_dma_mm_read_address
	wire          dma_fifo_subsystem_3_dma_mm_read_read;                                   // dma_fifo_subsystem_3:dma_mm_read_read -> mm_interconnect_0:dma_fifo_subsystem_3_dma_mm_read_read
	wire   [31:0] dma_fifo_subsystem_3_dma_mm_read_byteenable;                             // dma_fifo_subsystem_3:dma_mm_read_byteenable -> mm_interconnect_0:dma_fifo_subsystem_3_dma_mm_read_byteenable
	wire          dma_fifo_subsystem_3_dma_mm_read_readdatavalid;                          // mm_interconnect_0:dma_fifo_subsystem_3_dma_mm_read_readdatavalid -> dma_fifo_subsystem_3:dma_mm_read_readdatavalid
	wire   [10:0] dma_fifo_subsystem_3_dma_mm_read_burstcount;                             // dma_fifo_subsystem_3:dma_mm_read_burstcount -> mm_interconnect_0:dma_fifo_subsystem_3_dma_mm_read_burstcount
	wire          mm_interconnect_0_ddr2_ram_avl_beginbursttransfer;                       // mm_interconnect_0:ddr2_ram_avl_beginbursttransfer -> ddr2_ram:avl_burstbegin
	wire  [255:0] mm_interconnect_0_ddr2_ram_avl_readdata;                                 // ddr2_ram:avl_rdata -> mm_interconnect_0:ddr2_ram_avl_readdata
	wire          mm_interconnect_0_ddr2_ram_avl_waitrequest;                              // ddr2_ram:avl_ready -> mm_interconnect_0:ddr2_ram_avl_waitrequest
	wire   [24:0] mm_interconnect_0_ddr2_ram_avl_address;                                  // mm_interconnect_0:ddr2_ram_avl_address -> ddr2_ram:avl_addr
	wire          mm_interconnect_0_ddr2_ram_avl_read;                                     // mm_interconnect_0:ddr2_ram_avl_read -> ddr2_ram:avl_read_req
	wire   [31:0] mm_interconnect_0_ddr2_ram_avl_byteenable;                               // mm_interconnect_0:ddr2_ram_avl_byteenable -> ddr2_ram:avl_be
	wire          mm_interconnect_0_ddr2_ram_avl_readdatavalid;                            // ddr2_ram:avl_rdata_valid -> mm_interconnect_0:ddr2_ram_avl_readdatavalid
	wire          mm_interconnect_0_ddr2_ram_avl_write;                                    // mm_interconnect_0:ddr2_ram_avl_write -> ddr2_ram:avl_write_req
	wire  [255:0] mm_interconnect_0_ddr2_ram_avl_writedata;                                // mm_interconnect_0:ddr2_ram_avl_writedata -> ddr2_ram:avl_wdata
	wire    [2:0] mm_interconnect_0_ddr2_ram_avl_burstcount;                               // mm_interconnect_0:ddr2_ram_avl_burstcount -> ddr2_ram:avl_size
	wire          mm_interconnect_0_ddr2_ram_1_avl_beginbursttransfer;                     // mm_interconnect_0:ddr2_ram_1_avl_beginbursttransfer -> ddr2_ram_1:avl_burstbegin
	wire  [255:0] mm_interconnect_0_ddr2_ram_1_avl_readdata;                               // ddr2_ram_1:avl_rdata -> mm_interconnect_0:ddr2_ram_1_avl_readdata
	wire          mm_interconnect_0_ddr2_ram_1_avl_waitrequest;                            // ddr2_ram_1:avl_ready -> mm_interconnect_0:ddr2_ram_1_avl_waitrequest
	wire   [24:0] mm_interconnect_0_ddr2_ram_1_avl_address;                                // mm_interconnect_0:ddr2_ram_1_avl_address -> ddr2_ram_1:avl_addr
	wire          mm_interconnect_0_ddr2_ram_1_avl_read;                                   // mm_interconnect_0:ddr2_ram_1_avl_read -> ddr2_ram_1:avl_read_req
	wire   [31:0] mm_interconnect_0_ddr2_ram_1_avl_byteenable;                             // mm_interconnect_0:ddr2_ram_1_avl_byteenable -> ddr2_ram_1:avl_be
	wire          mm_interconnect_0_ddr2_ram_1_avl_readdatavalid;                          // ddr2_ram_1:avl_rdata_valid -> mm_interconnect_0:ddr2_ram_1_avl_readdatavalid
	wire          mm_interconnect_0_ddr2_ram_1_avl_write;                                  // mm_interconnect_0:ddr2_ram_1_avl_write -> ddr2_ram_1:avl_write_req
	wire  [255:0] mm_interconnect_0_ddr2_ram_1_avl_writedata;                              // mm_interconnect_0:ddr2_ram_1_avl_writedata -> ddr2_ram_1:avl_wdata
	wire    [2:0] mm_interconnect_0_ddr2_ram_1_avl_burstcount;                             // mm_interconnect_0:ddr2_ram_1_avl_burstcount -> ddr2_ram_1:avl_size
	wire          ddr2_ram_1_afi_clk_clk;                                                  // ddr2_ram_1:afi_clk -> [mm_interconnect_0:ddr2_ram_1_afi_clk_clk, rst_controller_003:clk]
	wire   [31:0] mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_readdata;                  // from_ETH_to_DDR:ETH_DMA_csr_readdata -> mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_csr_readdata
	wire    [2:0] mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_address;                   // mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_csr_address -> from_ETH_to_DDR:ETH_DMA_csr_address
	wire          mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_read;                      // mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_csr_read -> from_ETH_to_DDR:ETH_DMA_csr_read
	wire    [3:0] mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_byteenable;                // mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_csr_byteenable -> from_ETH_to_DDR:ETH_DMA_csr_byteenable
	wire          mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_write;                     // mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_csr_write -> from_ETH_to_DDR:ETH_DMA_csr_write
	wire   [31:0] mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_writedata;                 // mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_csr_writedata -> from_ETH_to_DDR:ETH_DMA_csr_writedata
	wire          mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_waitrequest;  // from_ETH_to_DDR:ETH_DMA_descriptor_slave_waitrequest -> mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_byteenable;   // mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_descriptor_slave_byteenable -> from_ETH_to_DDR:ETH_DMA_descriptor_slave_byteenable
	wire          mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_write;        // mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_descriptor_slave_write -> from_ETH_to_DDR:ETH_DMA_descriptor_slave_write
	wire  [127:0] mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_writedata;    // mm_interconnect_0:from_ETH_to_DDR_ETH_DMA_descriptor_slave_writedata -> from_ETH_to_DDR:ETH_DMA_descriptor_slave_writedata
	wire          mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                     // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                       // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                    // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                        // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire          mm_interconnect_0_jtag_avalon_jtag_slave_read;                           // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire          mm_interconnect_0_jtag_avalon_jtag_slave_write;                          // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                      // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire   [31:0] mm_interconnect_0_nios_cpu_debug_mem_slave_readdata;                     // nios_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios_cpu_debug_mem_slave_readdata
	wire          mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest;                  // nios_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_cpu_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess;                  // mm_interconnect_0:nios_cpu_debug_mem_slave_debugaccess -> nios_cpu:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_nios_cpu_debug_mem_slave_address;                      // mm_interconnect_0:nios_cpu_debug_mem_slave_address -> nios_cpu:debug_mem_slave_address
	wire          mm_interconnect_0_nios_cpu_debug_mem_slave_read;                         // mm_interconnect_0:nios_cpu_debug_mem_slave_read -> nios_cpu:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable;                   // mm_interconnect_0:nios_cpu_debug_mem_slave_byteenable -> nios_cpu:debug_mem_slave_byteenable
	wire          mm_interconnect_0_nios_cpu_debug_mem_slave_write;                        // mm_interconnect_0:nios_cpu_debug_mem_slave_write -> nios_cpu:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_nios_cpu_debug_mem_slave_writedata;                    // mm_interconnect_0:nios_cpu_debug_mem_slave_writedata -> nios_cpu:debug_mem_slave_writedata
	wire   [31:0] mm_interconnect_0_dma_fifo_susbystem_dma_csr_readdata;                   // dma_fifo_susbystem:dma_csr_readdata -> mm_interconnect_0:dma_fifo_susbystem_dma_csr_readdata
	wire    [2:0] mm_interconnect_0_dma_fifo_susbystem_dma_csr_address;                    // mm_interconnect_0:dma_fifo_susbystem_dma_csr_address -> dma_fifo_susbystem:dma_csr_address
	wire          mm_interconnect_0_dma_fifo_susbystem_dma_csr_read;                       // mm_interconnect_0:dma_fifo_susbystem_dma_csr_read -> dma_fifo_susbystem:dma_csr_read
	wire    [3:0] mm_interconnect_0_dma_fifo_susbystem_dma_csr_byteenable;                 // mm_interconnect_0:dma_fifo_susbystem_dma_csr_byteenable -> dma_fifo_susbystem:dma_csr_byteenable
	wire          mm_interconnect_0_dma_fifo_susbystem_dma_csr_write;                      // mm_interconnect_0:dma_fifo_susbystem_dma_csr_write -> dma_fifo_susbystem:dma_csr_write
	wire   [31:0] mm_interconnect_0_dma_fifo_susbystem_dma_csr_writedata;                  // mm_interconnect_0:dma_fifo_susbystem_dma_csr_writedata -> dma_fifo_susbystem:dma_csr_writedata
	wire   [31:0] mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_readdata;                 // dma_fifo_subsystem_1:dma_csr_readdata -> mm_interconnect_0:dma_fifo_subsystem_1_dma_csr_readdata
	wire    [2:0] mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_address;                  // mm_interconnect_0:dma_fifo_subsystem_1_dma_csr_address -> dma_fifo_subsystem_1:dma_csr_address
	wire          mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_read;                     // mm_interconnect_0:dma_fifo_subsystem_1_dma_csr_read -> dma_fifo_subsystem_1:dma_csr_read
	wire    [3:0] mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_byteenable;               // mm_interconnect_0:dma_fifo_subsystem_1_dma_csr_byteenable -> dma_fifo_subsystem_1:dma_csr_byteenable
	wire          mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_write;                    // mm_interconnect_0:dma_fifo_subsystem_1_dma_csr_write -> dma_fifo_subsystem_1:dma_csr_write
	wire   [31:0] mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_writedata;                // mm_interconnect_0:dma_fifo_subsystem_1_dma_csr_writedata -> dma_fifo_subsystem_1:dma_csr_writedata
	wire   [31:0] mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_readdata;                 // dma_fifo_subsystem_2:dma_csr_readdata -> mm_interconnect_0:dma_fifo_subsystem_2_dma_csr_readdata
	wire    [2:0] mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_address;                  // mm_interconnect_0:dma_fifo_subsystem_2_dma_csr_address -> dma_fifo_subsystem_2:dma_csr_address
	wire          mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_read;                     // mm_interconnect_0:dma_fifo_subsystem_2_dma_csr_read -> dma_fifo_subsystem_2:dma_csr_read
	wire    [3:0] mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_byteenable;               // mm_interconnect_0:dma_fifo_subsystem_2_dma_csr_byteenable -> dma_fifo_subsystem_2:dma_csr_byteenable
	wire          mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_write;                    // mm_interconnect_0:dma_fifo_subsystem_2_dma_csr_write -> dma_fifo_subsystem_2:dma_csr_write
	wire   [31:0] mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_writedata;                // mm_interconnect_0:dma_fifo_subsystem_2_dma_csr_writedata -> dma_fifo_subsystem_2:dma_csr_writedata
	wire   [31:0] mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_readdata;                 // dma_fifo_subsystem_3:dma_csr_readdata -> mm_interconnect_0:dma_fifo_subsystem_3_dma_csr_readdata
	wire    [2:0] mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_address;                  // mm_interconnect_0:dma_fifo_subsystem_3_dma_csr_address -> dma_fifo_subsystem_3:dma_csr_address
	wire          mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_read;                     // mm_interconnect_0:dma_fifo_subsystem_3_dma_csr_read -> dma_fifo_subsystem_3:dma_csr_read
	wire    [3:0] mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_byteenable;               // mm_interconnect_0:dma_fifo_subsystem_3_dma_csr_byteenable -> dma_fifo_subsystem_3:dma_csr_byteenable
	wire          mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_write;                    // mm_interconnect_0:dma_fifo_subsystem_3_dma_csr_write -> dma_fifo_subsystem_3:dma_csr_write
	wire   [31:0] mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_writedata;                // mm_interconnect_0:dma_fifo_subsystem_3_dma_csr_writedata -> dma_fifo_subsystem_3:dma_csr_writedata
	wire   [31:0] mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_readdata;                 // dma_fifo_subsystem_4:dma_csr_readdata -> mm_interconnect_0:dma_fifo_subsystem_4_dma_csr_readdata
	wire    [2:0] mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_address;                  // mm_interconnect_0:dma_fifo_subsystem_4_dma_csr_address -> dma_fifo_subsystem_4:dma_csr_address
	wire          mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_read;                     // mm_interconnect_0:dma_fifo_subsystem_4_dma_csr_read -> dma_fifo_subsystem_4:dma_csr_read
	wire    [3:0] mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_byteenable;               // mm_interconnect_0:dma_fifo_subsystem_4_dma_csr_byteenable -> dma_fifo_subsystem_4:dma_csr_byteenable
	wire          mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_write;                    // mm_interconnect_0:dma_fifo_subsystem_4_dma_csr_write -> dma_fifo_subsystem_4:dma_csr_write
	wire   [31:0] mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_writedata;                // mm_interconnect_0:dma_fifo_subsystem_4_dma_csr_writedata -> dma_fifo_subsystem_4:dma_csr_writedata
	wire          mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_waitrequest;   // dma_fifo_susbystem:dma_descriptor_slave_waitrequest -> mm_interconnect_0:dma_fifo_susbystem_dma_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_byteenable;    // mm_interconnect_0:dma_fifo_susbystem_dma_descriptor_slave_byteenable -> dma_fifo_susbystem:dma_descriptor_slave_byteenable
	wire          mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_write;         // mm_interconnect_0:dma_fifo_susbystem_dma_descriptor_slave_write -> dma_fifo_susbystem:dma_descriptor_slave_write
	wire  [127:0] mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_writedata;     // mm_interconnect_0:dma_fifo_susbystem_dma_descriptor_slave_writedata -> dma_fifo_susbystem:dma_descriptor_slave_writedata
	wire          mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_waitrequest; // dma_fifo_subsystem_1:dma_descriptor_slave_waitrequest -> mm_interconnect_0:dma_fifo_subsystem_1_dma_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_byteenable;  // mm_interconnect_0:dma_fifo_subsystem_1_dma_descriptor_slave_byteenable -> dma_fifo_subsystem_1:dma_descriptor_slave_byteenable
	wire          mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_write;       // mm_interconnect_0:dma_fifo_subsystem_1_dma_descriptor_slave_write -> dma_fifo_subsystem_1:dma_descriptor_slave_write
	wire  [127:0] mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_writedata;   // mm_interconnect_0:dma_fifo_subsystem_1_dma_descriptor_slave_writedata -> dma_fifo_subsystem_1:dma_descriptor_slave_writedata
	wire          mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_waitrequest; // dma_fifo_subsystem_2:dma_descriptor_slave_waitrequest -> mm_interconnect_0:dma_fifo_subsystem_2_dma_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_byteenable;  // mm_interconnect_0:dma_fifo_subsystem_2_dma_descriptor_slave_byteenable -> dma_fifo_subsystem_2:dma_descriptor_slave_byteenable
	wire          mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_write;       // mm_interconnect_0:dma_fifo_subsystem_2_dma_descriptor_slave_write -> dma_fifo_subsystem_2:dma_descriptor_slave_write
	wire  [127:0] mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_writedata;   // mm_interconnect_0:dma_fifo_subsystem_2_dma_descriptor_slave_writedata -> dma_fifo_subsystem_2:dma_descriptor_slave_writedata
	wire          mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_waitrequest; // dma_fifo_subsystem_3:dma_descriptor_slave_waitrequest -> mm_interconnect_0:dma_fifo_subsystem_3_dma_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_byteenable;  // mm_interconnect_0:dma_fifo_subsystem_3_dma_descriptor_slave_byteenable -> dma_fifo_subsystem_3:dma_descriptor_slave_byteenable
	wire          mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_write;       // mm_interconnect_0:dma_fifo_subsystem_3_dma_descriptor_slave_write -> dma_fifo_subsystem_3:dma_descriptor_slave_write
	wire  [127:0] mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_writedata;   // mm_interconnect_0:dma_fifo_subsystem_3_dma_descriptor_slave_writedata -> dma_fifo_subsystem_3:dma_descriptor_slave_writedata
	wire          mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_waitrequest; // dma_fifo_subsystem_4:dma_descriptor_slave_waitrequest -> mm_interconnect_0:dma_fifo_subsystem_4_dma_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_byteenable;  // mm_interconnect_0:dma_fifo_subsystem_4_dma_descriptor_slave_byteenable -> dma_fifo_subsystem_4:dma_descriptor_slave_byteenable
	wire          mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_write;       // mm_interconnect_0:dma_fifo_subsystem_4_dma_descriptor_slave_write -> dma_fifo_subsystem_4:dma_descriptor_slave_write
	wire  [127:0] mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_writedata;   // mm_interconnect_0:dma_fifo_subsystem_4_dma_descriptor_slave_writedata -> dma_fifo_subsystem_4:dma_descriptor_slave_writedata
	wire          mm_interconnect_0_system_ram_s1_chipselect;                              // mm_interconnect_0:system_ram_s1_chipselect -> system_ram:chipselect
	wire   [31:0] mm_interconnect_0_system_ram_s1_readdata;                                // system_ram:readdata -> mm_interconnect_0:system_ram_s1_readdata
	wire   [16:0] mm_interconnect_0_system_ram_s1_address;                                 // mm_interconnect_0:system_ram_s1_address -> system_ram:address
	wire    [3:0] mm_interconnect_0_system_ram_s1_byteenable;                              // mm_interconnect_0:system_ram_s1_byteenable -> system_ram:byteenable
	wire          mm_interconnect_0_system_ram_s1_write;                                   // mm_interconnect_0:system_ram_s1_write -> system_ram:write
	wire   [31:0] mm_interconnect_0_system_ram_s1_writedata;                               // mm_interconnect_0:system_ram_s1_writedata -> system_ram:writedata
	wire          mm_interconnect_0_system_ram_s1_clken;                                   // mm_interconnect_0:system_ram_s1_clken -> system_ram:clken
	wire          mm_interconnect_0_ctrl_sig_s1_chipselect;                                // mm_interconnect_0:ctrl_sig_s1_chipselect -> ctrl_sig:chipselect
	wire   [31:0] mm_interconnect_0_ctrl_sig_s1_readdata;                                  // ctrl_sig:readdata -> mm_interconnect_0:ctrl_sig_s1_readdata
	wire    [1:0] mm_interconnect_0_ctrl_sig_s1_address;                                   // mm_interconnect_0:ctrl_sig_s1_address -> ctrl_sig:address
	wire          mm_interconnect_0_ctrl_sig_s1_write;                                     // mm_interconnect_0:ctrl_sig_s1_write -> ctrl_sig:write_n
	wire   [31:0] mm_interconnect_0_ctrl_sig_s1_writedata;                                 // mm_interconnect_0:ctrl_sig_s1_writedata -> ctrl_sig:writedata
	wire          mm_interconnect_0_sys_timer_s1_chipselect;                               // mm_interconnect_0:sys_timer_s1_chipselect -> sys_timer:chipselect
	wire   [15:0] mm_interconnect_0_sys_timer_s1_readdata;                                 // sys_timer:readdata -> mm_interconnect_0:sys_timer_s1_readdata
	wire    [2:0] mm_interconnect_0_sys_timer_s1_address;                                  // mm_interconnect_0:sys_timer_s1_address -> sys_timer:address
	wire          mm_interconnect_0_sys_timer_s1_write;                                    // mm_interconnect_0:sys_timer_s1_write -> sys_timer:write_n
	wire   [15:0] mm_interconnect_0_sys_timer_s1_writedata;                                // mm_interconnect_0:sys_timer_s1_writedata -> sys_timer:writedata
	wire          mm_interconnect_0_pilot_sig_s1_chipselect;                               // mm_interconnect_0:pilot_sig_s1_chipselect -> pilot_sig:chipselect
	wire   [31:0] mm_interconnect_0_pilot_sig_s1_readdata;                                 // pilot_sig:readdata -> mm_interconnect_0:pilot_sig_s1_readdata
	wire    [1:0] mm_interconnect_0_pilot_sig_s1_address;                                  // mm_interconnect_0:pilot_sig_s1_address -> pilot_sig:address
	wire          mm_interconnect_0_pilot_sig_s1_write;                                    // mm_interconnect_0:pilot_sig_s1_write -> pilot_sig:write_n
	wire   [31:0] mm_interconnect_0_pilot_sig_s1_writedata;                                // mm_interconnect_0:pilot_sig_s1_writedata -> pilot_sig:writedata
	wire          mm_interconnect_0_input_io_s1_chipselect;                                // mm_interconnect_0:input_IO_s1_chipselect -> input_IO:chipselect
	wire   [31:0] mm_interconnect_0_input_io_s1_readdata;                                  // input_IO:readdata -> mm_interconnect_0:input_IO_s1_readdata
	wire    [1:0] mm_interconnect_0_input_io_s1_address;                                   // mm_interconnect_0:input_IO_s1_address -> input_IO:address
	wire          mm_interconnect_0_input_io_s1_write;                                     // mm_interconnect_0:input_IO_s1_write -> input_IO:write_n
	wire   [31:0] mm_interconnect_0_input_io_s1_writedata;                                 // mm_interconnect_0:input_IO_s1_writedata -> input_IO:writedata
	wire          mm_interconnect_0_input_io_0_s1_chipselect;                              // mm_interconnect_0:input_IO_0_s1_chipselect -> input_IO_0:chipselect
	wire   [31:0] mm_interconnect_0_input_io_0_s1_readdata;                                // input_IO_0:readdata -> mm_interconnect_0:input_IO_0_s1_readdata
	wire    [1:0] mm_interconnect_0_input_io_0_s1_address;                                 // mm_interconnect_0:input_IO_0_s1_address -> input_IO_0:address
	wire          mm_interconnect_0_input_io_0_s1_write;                                   // mm_interconnect_0:input_IO_0_s1_write -> input_IO_0:write_n
	wire   [31:0] mm_interconnect_0_input_io_0_s1_writedata;                               // mm_interconnect_0:input_IO_0_s1_writedata -> input_IO_0:writedata
	wire          mm_interconnect_0_input_io_1_s1_chipselect;                              // mm_interconnect_0:input_IO_1_s1_chipselect -> input_IO_1:chipselect
	wire   [31:0] mm_interconnect_0_input_io_1_s1_readdata;                                // input_IO_1:readdata -> mm_interconnect_0:input_IO_1_s1_readdata
	wire    [1:0] mm_interconnect_0_input_io_1_s1_address;                                 // mm_interconnect_0:input_IO_1_s1_address -> input_IO_1:address
	wire          mm_interconnect_0_input_io_1_s1_write;                                   // mm_interconnect_0:input_IO_1_s1_write -> input_IO_1:write_n
	wire   [31:0] mm_interconnect_0_input_io_1_s1_writedata;                               // mm_interconnect_0:input_IO_1_s1_writedata -> input_IO_1:writedata
	wire          mm_interconnect_0_input_io_2_s1_chipselect;                              // mm_interconnect_0:input_IO_2_s1_chipselect -> input_IO_2:chipselect
	wire   [31:0] mm_interconnect_0_input_io_2_s1_readdata;                                // input_IO_2:readdata -> mm_interconnect_0:input_IO_2_s1_readdata
	wire    [1:0] mm_interconnect_0_input_io_2_s1_address;                                 // mm_interconnect_0:input_IO_2_s1_address -> input_IO_2:address
	wire          mm_interconnect_0_input_io_2_s1_write;                                   // mm_interconnect_0:input_IO_2_s1_write -> input_IO_2:write_n
	wire   [31:0] mm_interconnect_0_input_io_2_s1_writedata;                               // mm_interconnect_0:input_IO_2_s1_writedata -> input_IO_2:writedata
	wire          mm_interconnect_0_input_io_3_s1_chipselect;                              // mm_interconnect_0:input_IO_3_s1_chipselect -> input_IO_3:chipselect
	wire   [31:0] mm_interconnect_0_input_io_3_s1_readdata;                                // input_IO_3:readdata -> mm_interconnect_0:input_IO_3_s1_readdata
	wire    [1:0] mm_interconnect_0_input_io_3_s1_address;                                 // mm_interconnect_0:input_IO_3_s1_address -> input_IO_3:address
	wire          mm_interconnect_0_input_io_3_s1_write;                                   // mm_interconnect_0:input_IO_3_s1_write -> input_IO_3:write_n
	wire   [31:0] mm_interconnect_0_input_io_3_s1_writedata;                               // mm_interconnect_0:input_IO_3_s1_writedata -> input_IO_3:writedata
	wire          mm_interconnect_0_input_io_4_s1_chipselect;                              // mm_interconnect_0:input_IO_4_s1_chipselect -> input_IO_4:chipselect
	wire   [31:0] mm_interconnect_0_input_io_4_s1_readdata;                                // input_IO_4:readdata -> mm_interconnect_0:input_IO_4_s1_readdata
	wire    [1:0] mm_interconnect_0_input_io_4_s1_address;                                 // mm_interconnect_0:input_IO_4_s1_address -> input_IO_4:address
	wire          mm_interconnect_0_input_io_4_s1_write;                                   // mm_interconnect_0:input_IO_4_s1_write -> input_IO_4:write_n
	wire   [31:0] mm_interconnect_0_input_io_4_s1_writedata;                               // mm_interconnect_0:input_IO_4_s1_writedata -> input_IO_4:writedata
	wire          mm_interconnect_0_input_io_5_s1_chipselect;                              // mm_interconnect_0:input_IO_5_s1_chipselect -> input_IO_5:chipselect
	wire   [31:0] mm_interconnect_0_input_io_5_s1_readdata;                                // input_IO_5:readdata -> mm_interconnect_0:input_IO_5_s1_readdata
	wire    [1:0] mm_interconnect_0_input_io_5_s1_address;                                 // mm_interconnect_0:input_IO_5_s1_address -> input_IO_5:address
	wire          mm_interconnect_0_input_io_5_s1_write;                                   // mm_interconnect_0:input_IO_5_s1_write -> input_IO_5:write_n
	wire   [31:0] mm_interconnect_0_input_io_5_s1_writedata;                               // mm_interconnect_0:input_IO_5_s1_writedata -> input_IO_5:writedata
	wire          irq_mapper_receiver0_irq;                                                // from_ETH_to_DDR:ETH_DMA_csr_irq_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                // dma_fifo_susbystem:dma_csr_irq_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                // dma_fifo_subsystem_1:dma_csr_irq_irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                // dma_fifo_subsystem_2:dma_csr_irq_irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                // dma_fifo_subsystem_3:dma_csr_irq_irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                // dma_fifo_subsystem_4:dma_csr_irq_irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                // jtag:av_irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver7_irq;                                                // sys_timer:irq -> irq_mapper:receiver7_irq
	wire          irq_mapper_receiver8_irq;                                                // pilot_sig:irq -> irq_mapper:receiver8_irq
	wire   [31:0] nios_cpu_irq_irq;                                                        // irq_mapper:sender_irq -> nios_cpu:irq
	wire          rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [ctrl_sig:reset_n, dma_fifo_subsystem_1:dma_reset_n_reset_n, dma_fifo_subsystem_1:fifo_stream_reset_reset_n, dma_fifo_subsystem_2:dma_reset_n_reset_n, dma_fifo_subsystem_2:fifo_stream_reset_reset_n, dma_fifo_subsystem_3:dma_reset_n_reset_n, dma_fifo_subsystem_3:fifo_stream_reset_reset_n, dma_fifo_subsystem_4:dma_reset_n_reset_n, dma_fifo_subsystem_4:fifo_stream_reset_reset_n, dma_fifo_susbystem:dma_reset_n_reset_n, dma_fifo_susbystem:fifo_stream_reset_reset_n, input_IO:reset_n, input_IO_0:reset_n, input_IO_1:reset_n, input_IO_2:reset_n, input_IO_3:reset_n, input_IO_4:reset_n, input_IO_5:reset_n, irq_mapper:reset, jtag:rst_n, mm_interconnect_0:from_ETH_to_DDR_reset_reset_bridge_in_reset_reset, mm_interconnect_0:nios_cpu_reset_reset_bridge_in_reset_reset, nios_cpu:reset_n, pilot_sig:reset_n, rst_translator:in_reset, sys_timer:reset_n, system_ram:reset]
	wire          rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [nios_cpu:reset_req, rst_translator:reset_req_in, system_ram:reset_req]
	wire          rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> ddr2_ram:soft_reset_n
	wire          nios_cpu_debug_reset_request_reset;                                      // nios_cpu:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1]
	wire          rst_controller_002_reset_out_reset;                                      // rst_controller_002:reset_out -> ddr2_ram_1:soft_reset_n
	wire          rst_controller_003_reset_out_reset;                                      // rst_controller_003:reset_out -> [mm_interconnect_0:ddr2_ram_1_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:ddr2_ram_1_soft_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_004_reset_out_reset;                                      // rst_controller_004:reset_out -> [mm_interconnect_0:ddr2_ram_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:ddr2_ram_soft_reset_reset_bridge_in_reset_reset]

	testbench_ls_ctrl_sig ctrl_sig (
		.clk        (clk_200_out_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_ctrl_sig_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ctrl_sig_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ctrl_sig_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ctrl_sig_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ctrl_sig_s1_readdata),   //                    .readdata
		.out_port   (ctrl_sig_export)                           // external_connection.export
	);

	testbench_ls_ddr2_ram ddr2_ram (
		.pll_ref_clk        (clk_50_clk),                                        //      pll_ref_clk.clk
		.global_reset_n     (reset_reset_n),                                     //     global_reset.reset_n
		.soft_reset_n       (~rst_controller_001_reset_out_reset),               //       soft_reset.reset_n
		.afi_clk            (clk_200_out_clk_clk),                               //          afi_clk.clk
		.afi_half_clk       (),                                                  //     afi_half_clk.clk
		.afi_reset_n        (),                                                  //        afi_reset.reset_n
		.afi_reset_export_n (),                                                  // afi_reset_export.reset_n
		.mem_a              (memory_mem_a),                                      //           memory.mem_a
		.mem_ba             (memory_mem_ba),                                     //                 .mem_ba
		.mem_ck             (memory_mem_ck),                                     //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                                   //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),                                    //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                                   //                 .mem_cs_n
		.mem_dm             (memory_mem_dm),                                     //                 .mem_dm
		.mem_ras_n          (memory_mem_ras_n),                                  //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                                  //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                                   //                 .mem_we_n
		.mem_dq             (memory_mem_dq),                                     //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),                                    //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                                  //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),                                    //                 .mem_odt
		.avl_ready          (mm_interconnect_0_ddr2_ram_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (mm_interconnect_0_ddr2_ram_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (mm_interconnect_0_ddr2_ram_avl_address),            //                 .address
		.avl_rdata_valid    (mm_interconnect_0_ddr2_ram_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (mm_interconnect_0_ddr2_ram_avl_readdata),           //                 .readdata
		.avl_wdata          (mm_interconnect_0_ddr2_ram_avl_writedata),          //                 .writedata
		.avl_be             (mm_interconnect_0_ddr2_ram_avl_byteenable),         //                 .byteenable
		.avl_read_req       (mm_interconnect_0_ddr2_ram_avl_read),               //                 .read
		.avl_write_req      (mm_interconnect_0_ddr2_ram_avl_write),              //                 .write
		.avl_size           (mm_interconnect_0_ddr2_ram_avl_burstcount),         //                 .burstcount
		.local_init_done    (ddr2_ram_status_local_init_done),                   //           status.local_init_done
		.local_cal_success  (ddr2_ram_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail     (ddr2_ram_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rdn            (oct_rdn),                                           //              oct.rdn
		.oct_rup            (oct_rup)                                            //                 .rup
	);

	testbench_ls_ddr2_ram ddr2_ram_1 (
		.pll_ref_clk        (clk_50_clk),                                          //      pll_ref_clk.clk
		.global_reset_n     (reset_reset_n),                                       //     global_reset.reset_n
		.soft_reset_n       (~rst_controller_002_reset_out_reset),                 //       soft_reset.reset_n
		.afi_clk            (ddr2_ram_1_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk       (),                                                    //     afi_half_clk.clk
		.afi_reset_n        (),                                                    //        afi_reset.reset_n
		.afi_reset_export_n (),                                                    // afi_reset_export.reset_n
		.mem_a              (memory_1_mem_a),                                      //           memory.mem_a
		.mem_ba             (memory_1_mem_ba),                                     //                 .mem_ba
		.mem_ck             (memory_1_mem_ck),                                     //                 .mem_ck
		.mem_ck_n           (memory_1_mem_ck_n),                                   //                 .mem_ck_n
		.mem_cke            (memory_1_mem_cke),                                    //                 .mem_cke
		.mem_cs_n           (memory_1_mem_cs_n),                                   //                 .mem_cs_n
		.mem_dm             (memory_1_mem_dm),                                     //                 .mem_dm
		.mem_ras_n          (memory_1_mem_ras_n),                                  //                 .mem_ras_n
		.mem_cas_n          (memory_1_mem_cas_n),                                  //                 .mem_cas_n
		.mem_we_n           (memory_1_mem_we_n),                                   //                 .mem_we_n
		.mem_dq             (memory_1_mem_dq),                                     //                 .mem_dq
		.mem_dqs            (memory_1_mem_dqs),                                    //                 .mem_dqs
		.mem_dqs_n          (memory_1_mem_dqs_n),                                  //                 .mem_dqs_n
		.mem_odt            (memory_1_mem_odt),                                    //                 .mem_odt
		.avl_ready          (mm_interconnect_0_ddr2_ram_1_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (mm_interconnect_0_ddr2_ram_1_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (mm_interconnect_0_ddr2_ram_1_avl_address),            //                 .address
		.avl_rdata_valid    (mm_interconnect_0_ddr2_ram_1_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (mm_interconnect_0_ddr2_ram_1_avl_readdata),           //                 .readdata
		.avl_wdata          (mm_interconnect_0_ddr2_ram_1_avl_writedata),          //                 .writedata
		.avl_be             (mm_interconnect_0_ddr2_ram_1_avl_byteenable),         //                 .byteenable
		.avl_read_req       (mm_interconnect_0_ddr2_ram_1_avl_read),               //                 .read
		.avl_write_req      (mm_interconnect_0_ddr2_ram_1_avl_write),              //                 .write
		.avl_size           (mm_interconnect_0_ddr2_ram_1_avl_burstcount),         //                 .burstcount
		.local_init_done    (),                                                    //           status.local_init_done
		.local_cal_success  (),                                                    //                 .local_cal_success
		.local_cal_fail     (),                                                    //                 .local_cal_fail
		.oct_rdn            (oct_1_rdn),                                           //              oct.rdn
		.oct_rup            (oct_1_rup)                                            //                 .rup
	);

	testbench_ls_dma_fifo_subsystem_1 dma_fifo_subsystem_1 (
		.dma_clock_clk                      (clk_200_out_clk_clk),                                                     //               dma_clock.clk
		.dma_csr_writedata                  (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_writedata),                //                 dma_csr.writedata
		.dma_csr_write                      (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_write),                    //                        .write
		.dma_csr_byteenable                 (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_byteenable),               //                        .byteenable
		.dma_csr_readdata                   (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_readdata),                 //                        .readdata
		.dma_csr_read                       (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_read),                     //                        .read
		.dma_csr_address                    (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_address),                  //                        .address
		.dma_csr_irq_irq                    (irq_mapper_receiver2_irq),                                                //             dma_csr_irq.irq
		.dma_descriptor_slave_write         (mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_write),       //    dma_descriptor_slave.write
		.dma_descriptor_slave_waitrequest   (mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_waitrequest), //                        .waitrequest
		.dma_descriptor_slave_writedata     (mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_writedata),   //                        .writedata
		.dma_descriptor_slave_byteenable    (mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_byteenable),  //                        .byteenable
		.dma_mm_read_address                (dma_fifo_subsystem_1_dma_mm_read_address),                                //             dma_mm_read.address
		.dma_mm_read_read                   (dma_fifo_subsystem_1_dma_mm_read_read),                                   //                        .read
		.dma_mm_read_byteenable             (dma_fifo_subsystem_1_dma_mm_read_byteenable),                             //                        .byteenable
		.dma_mm_read_readdata               (dma_fifo_subsystem_1_dma_mm_read_readdata),                               //                        .readdata
		.dma_mm_read_waitrequest            (dma_fifo_subsystem_1_dma_mm_read_waitrequest),                            //                        .waitrequest
		.dma_mm_read_readdatavalid          (dma_fifo_subsystem_1_dma_mm_read_readdatavalid),                          //                        .readdatavalid
		.dma_mm_read_burstcount             (dma_fifo_subsystem_1_dma_mm_read_burstcount),                             //                        .burstcount
		.dma_reset_n_reset_n                (~rst_controller_reset_out_reset),                                         //             dma_reset_n.reset_n
		.fifo_stream_clock_clk              (clk_200_out_clk_clk),                                                     //       fifo_stream_clock.clk
		.fifo_stream_conduit_end_fifo_data  (fifo_stream_1_fifo_data),                                                 // fifo_stream_conduit_end.fifo_data
		.fifo_stream_conduit_end_fifo_write (fifo_stream_1_fifo_write),                                                //                        .fifo_write
		.fifo_stream_conduit_end_fifo_send  (fifo_stream_1_fifo_send),                                                 //                        .fifo_send
		.fifo_stream_reset_reset_n          (~rst_controller_reset_out_reset)                                          //       fifo_stream_reset.reset_n
	);

	testbench_ls_dma_fifo_subsystem_2 dma_fifo_subsystem_2 (
		.dma_clock_clk                      (clk_200_out_clk_clk),                                                     //               dma_clock.clk
		.dma_csr_writedata                  (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_writedata),                //                 dma_csr.writedata
		.dma_csr_write                      (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_write),                    //                        .write
		.dma_csr_byteenable                 (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_byteenable),               //                        .byteenable
		.dma_csr_readdata                   (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_readdata),                 //                        .readdata
		.dma_csr_read                       (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_read),                     //                        .read
		.dma_csr_address                    (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_address),                  //                        .address
		.dma_csr_irq_irq                    (irq_mapper_receiver3_irq),                                                //             dma_csr_irq.irq
		.dma_descriptor_slave_write         (mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_write),       //    dma_descriptor_slave.write
		.dma_descriptor_slave_waitrequest   (mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_waitrequest), //                        .waitrequest
		.dma_descriptor_slave_writedata     (mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_writedata),   //                        .writedata
		.dma_descriptor_slave_byteenable    (mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_byteenable),  //                        .byteenable
		.dma_mm_read_address                (dma_fifo_subsystem_2_dma_mm_read_address),                                //             dma_mm_read.address
		.dma_mm_read_read                   (dma_fifo_subsystem_2_dma_mm_read_read),                                   //                        .read
		.dma_mm_read_byteenable             (dma_fifo_subsystem_2_dma_mm_read_byteenable),                             //                        .byteenable
		.dma_mm_read_readdata               (dma_fifo_subsystem_2_dma_mm_read_readdata),                               //                        .readdata
		.dma_mm_read_waitrequest            (dma_fifo_subsystem_2_dma_mm_read_waitrequest),                            //                        .waitrequest
		.dma_mm_read_readdatavalid          (dma_fifo_subsystem_2_dma_mm_read_readdatavalid),                          //                        .readdatavalid
		.dma_mm_read_burstcount             (dma_fifo_subsystem_2_dma_mm_read_burstcount),                             //                        .burstcount
		.dma_reset_n_reset_n                (~rst_controller_reset_out_reset),                                         //             dma_reset_n.reset_n
		.fifo_stream_clock_clk              (clk_200_out_clk_clk),                                                     //       fifo_stream_clock.clk
		.fifo_stream_conduit_end_fifo_data  (dma_fifo_subsystem_2_fifo_stream_conduit_end_fifo_data),                  // fifo_stream_conduit_end.fifo_data
		.fifo_stream_conduit_end_fifo_write (dma_fifo_subsystem_2_fifo_stream_conduit_end_fifo_write),                 //                        .fifo_write
		.fifo_stream_conduit_end_fifo_send  (dma_fifo_subsystem_2_fifo_stream_conduit_end_fifo_send),                  //                        .fifo_send
		.fifo_stream_reset_reset_n          (~rst_controller_reset_out_reset)                                          //       fifo_stream_reset.reset_n
	);

	testbench_ls_dma_fifo_subsystem_3 dma_fifo_subsystem_3 (
		.dma_clock_clk                      (clk_200_out_clk_clk),                                                     //               dma_clock.clk
		.dma_csr_writedata                  (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_writedata),                //                 dma_csr.writedata
		.dma_csr_write                      (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_write),                    //                        .write
		.dma_csr_byteenable                 (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_byteenable),               //                        .byteenable
		.dma_csr_readdata                   (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_readdata),                 //                        .readdata
		.dma_csr_read                       (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_read),                     //                        .read
		.dma_csr_address                    (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_address),                  //                        .address
		.dma_csr_irq_irq                    (irq_mapper_receiver4_irq),                                                //             dma_csr_irq.irq
		.dma_descriptor_slave_write         (mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_write),       //    dma_descriptor_slave.write
		.dma_descriptor_slave_waitrequest   (mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_waitrequest), //                        .waitrequest
		.dma_descriptor_slave_writedata     (mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_writedata),   //                        .writedata
		.dma_descriptor_slave_byteenable    (mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_byteenable),  //                        .byteenable
		.dma_mm_read_address                (dma_fifo_subsystem_3_dma_mm_read_address),                                //             dma_mm_read.address
		.dma_mm_read_read                   (dma_fifo_subsystem_3_dma_mm_read_read),                                   //                        .read
		.dma_mm_read_byteenable             (dma_fifo_subsystem_3_dma_mm_read_byteenable),                             //                        .byteenable
		.dma_mm_read_readdata               (dma_fifo_subsystem_3_dma_mm_read_readdata),                               //                        .readdata
		.dma_mm_read_waitrequest            (dma_fifo_subsystem_3_dma_mm_read_waitrequest),                            //                        .waitrequest
		.dma_mm_read_readdatavalid          (dma_fifo_subsystem_3_dma_mm_read_readdatavalid),                          //                        .readdatavalid
		.dma_mm_read_burstcount             (dma_fifo_subsystem_3_dma_mm_read_burstcount),                             //                        .burstcount
		.dma_reset_n_reset_n                (~rst_controller_reset_out_reset),                                         //             dma_reset_n.reset_n
		.fifo_stream_clock_clk              (clk_200_out_clk_clk),                                                     //       fifo_stream_clock.clk
		.fifo_stream_conduit_end_fifo_data  (dma_fifo_subsystem_3_fifo_stream_conduit_end_fifo_data),                  // fifo_stream_conduit_end.fifo_data
		.fifo_stream_conduit_end_fifo_write (dma_fifo_subsystem_3_fifo_stream_conduit_end_fifo_write),                 //                        .fifo_write
		.fifo_stream_conduit_end_fifo_send  (dma_fifo_subsystem_3_fifo_stream_conduit_end_fifo_send),                  //                        .fifo_send
		.fifo_stream_reset_reset_n          (~rst_controller_reset_out_reset)                                          //       fifo_stream_reset.reset_n
	);

	testbench_ls_dma_fifo_subsystem_4 dma_fifo_subsystem_4 (
		.dma_clock_clk                      (clk_200_out_clk_clk),                                                     //               dma_clock.clk
		.dma_csr_writedata                  (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_writedata),                //                 dma_csr.writedata
		.dma_csr_write                      (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_write),                    //                        .write
		.dma_csr_byteenable                 (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_byteenable),               //                        .byteenable
		.dma_csr_readdata                   (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_readdata),                 //                        .readdata
		.dma_csr_read                       (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_read),                     //                        .read
		.dma_csr_address                    (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_address),                  //                        .address
		.dma_csr_irq_irq                    (irq_mapper_receiver5_irq),                                                //             dma_csr_irq.irq
		.dma_descriptor_slave_write         (mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_write),       //    dma_descriptor_slave.write
		.dma_descriptor_slave_waitrequest   (mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_waitrequest), //                        .waitrequest
		.dma_descriptor_slave_writedata     (mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_writedata),   //                        .writedata
		.dma_descriptor_slave_byteenable    (mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_byteenable),  //                        .byteenable
		.dma_mm_read_address                (dma_fifo_subsystem_4_dma_mm_read_address),                                //             dma_mm_read.address
		.dma_mm_read_read                   (dma_fifo_subsystem_4_dma_mm_read_read),                                   //                        .read
		.dma_mm_read_byteenable             (dma_fifo_subsystem_4_dma_mm_read_byteenable),                             //                        .byteenable
		.dma_mm_read_readdata               (dma_fifo_subsystem_4_dma_mm_read_readdata),                               //                        .readdata
		.dma_mm_read_waitrequest            (dma_fifo_subsystem_4_dma_mm_read_waitrequest),                            //                        .waitrequest
		.dma_mm_read_readdatavalid          (dma_fifo_subsystem_4_dma_mm_read_readdatavalid),                          //                        .readdatavalid
		.dma_mm_read_burstcount             (dma_fifo_subsystem_4_dma_mm_read_burstcount),                             //                        .burstcount
		.dma_reset_n_reset_n                (~rst_controller_reset_out_reset),                                         //             dma_reset_n.reset_n
		.fifo_stream_clock_clk              (clk_200_out_clk_clk),                                                     //       fifo_stream_clock.clk
		.fifo_stream_conduit_end_fifo_data  (dma_fifo_subsystem_4_fifo_stream_conduit_end_fifo_data),                  // fifo_stream_conduit_end.fifo_data
		.fifo_stream_conduit_end_fifo_write (dma_fifo_subsystem_4_fifo_stream_conduit_end_fifo_write),                 //                        .fifo_write
		.fifo_stream_conduit_end_fifo_send  (dma_fifo_subsystem_4_fifo_stream_conduit_end_fifo_send),                  //                        .fifo_send
		.fifo_stream_reset_reset_n          (~rst_controller_reset_out_reset)                                          //       fifo_stream_reset.reset_n
	);

	testbench_ls_dma_fifo_susbystem dma_fifo_susbystem (
		.dma_clock_clk                      (clk_200_out_clk_clk),                                                   //               dma_clock.clk
		.dma_csr_writedata                  (mm_interconnect_0_dma_fifo_susbystem_dma_csr_writedata),                //                 dma_csr.writedata
		.dma_csr_write                      (mm_interconnect_0_dma_fifo_susbystem_dma_csr_write),                    //                        .write
		.dma_csr_byteenable                 (mm_interconnect_0_dma_fifo_susbystem_dma_csr_byteenable),               //                        .byteenable
		.dma_csr_readdata                   (mm_interconnect_0_dma_fifo_susbystem_dma_csr_readdata),                 //                        .readdata
		.dma_csr_read                       (mm_interconnect_0_dma_fifo_susbystem_dma_csr_read),                     //                        .read
		.dma_csr_address                    (mm_interconnect_0_dma_fifo_susbystem_dma_csr_address),                  //                        .address
		.dma_csr_irq_irq                    (irq_mapper_receiver1_irq),                                              //             dma_csr_irq.irq
		.dma_descriptor_slave_write         (mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_write),       //    dma_descriptor_slave.write
		.dma_descriptor_slave_waitrequest   (mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_waitrequest), //                        .waitrequest
		.dma_descriptor_slave_writedata     (mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_writedata),   //                        .writedata
		.dma_descriptor_slave_byteenable    (mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_byteenable),  //                        .byteenable
		.dma_mm_read_address                (dma_fifo_susbystem_dma_mm_read_address),                                //             dma_mm_read.address
		.dma_mm_read_read                   (dma_fifo_susbystem_dma_mm_read_read),                                   //                        .read
		.dma_mm_read_byteenable             (dma_fifo_susbystem_dma_mm_read_byteenable),                             //                        .byteenable
		.dma_mm_read_readdata               (dma_fifo_susbystem_dma_mm_read_readdata),                               //                        .readdata
		.dma_mm_read_waitrequest            (dma_fifo_susbystem_dma_mm_read_waitrequest),                            //                        .waitrequest
		.dma_mm_read_readdatavalid          (dma_fifo_susbystem_dma_mm_read_readdatavalid),                          //                        .readdatavalid
		.dma_mm_read_burstcount             (dma_fifo_susbystem_dma_mm_read_burstcount),                             //                        .burstcount
		.dma_reset_n_reset_n                (~rst_controller_reset_out_reset),                                       //             dma_reset_n.reset_n
		.fifo_stream_clock_clk              (clk_200_out_clk_clk),                                                   //       fifo_stream_clock.clk
		.fifo_stream_conduit_end_fifo_data  (fifo_stream_fifo_data),                                                 // fifo_stream_conduit_end.fifo_data
		.fifo_stream_conduit_end_fifo_write (fifo_stream_fifo_write),                                                //                        .fifo_write
		.fifo_stream_conduit_end_fifo_send  (fifo_stream_fifo_send),                                                 //                        .fifo_send
		.fifo_stream_reset_reset_n          (~rst_controller_reset_out_reset)                                        //       fifo_stream_reset.reset_n
	);

	testbench_ls_from_ETH_to_DDR from_eth_to_ddr (
		.ETH_DMA_csr_writedata                (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_writedata),                //              ETH_DMA_csr.writedata
		.ETH_DMA_csr_write                    (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_write),                    //                         .write
		.ETH_DMA_csr_byteenable               (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_byteenable),               //                         .byteenable
		.ETH_DMA_csr_readdata                 (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_readdata),                 //                         .readdata
		.ETH_DMA_csr_read                     (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_read),                     //                         .read
		.ETH_DMA_csr_address                  (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_address),                  //                         .address
		.ETH_DMA_csr_irq_irq                  (irq_mapper_receiver0_irq),                                               //          ETH_DMA_csr_irq.irq
		.ETH_DMA_descriptor_slave_write       (mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_write),       // ETH_DMA_descriptor_slave.write
		.ETH_DMA_descriptor_slave_waitrequest (mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_waitrequest), //                         .waitrequest
		.ETH_DMA_descriptor_slave_writedata   (mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_writedata),   //                         .writedata
		.ETH_DMA_descriptor_slave_byteenable  (mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_byteenable),  //                         .byteenable
		.ETH_DMA_mm_write_address             (from_eth_to_ddr_eth_dma_mm_write_address),                               //         ETH_DMA_mm_write.address
		.ETH_DMA_mm_write_write               (from_eth_to_ddr_eth_dma_mm_write_write),                                 //                         .write
		.ETH_DMA_mm_write_byteenable          (from_eth_to_ddr_eth_dma_mm_write_byteenable),                            //                         .byteenable
		.ETH_DMA_mm_write_writedata           (from_eth_to_ddr_eth_dma_mm_write_writedata),                             //                         .writedata
		.ETH_DMA_mm_write_waitrequest         (from_eth_to_ddr_eth_dma_mm_write_waitrequest),                           //                         .waitrequest
		.clk_clk                              (clk_200_out_clk_clk),                                                    //                      clk.clk
		.eth_fifo_tofifo_fifo_data            (from_fifo_fifo_data),                                                    //          eth_fifo_tofifo.fifo_data
		.eth_fifo_tofifo_fifo_read            (from_fifo_fifo_read),                                                    //                         .fifo_read
		.eth_fifo_tofifo_fifo_empty           (from_fifo_fifo_empty),                                                   //                         .fifo_empty
		.eth_fifo_tofifo_fifo_full            (from_fifo_fifo_full),                                                    //                         .fifo_full
		.reset_reset_n                        (reset_reset_n)                                                           //                    reset.reset_n
	);

	testbench_ls_input_IO input_io (
		.clk        (clk_200_out_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_input_io_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_io_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_io_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_io_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_io_s1_readdata),   //                    .readdata
		.in_port    (input_io_external_connection_export)       // external_connection.export
	);

	testbench_ls_input_IO input_io_0 (
		.clk        (clk_200_out_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_input_io_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_io_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_io_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_io_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_io_0_s1_readdata),   //                    .readdata
		.in_port    (input_io_0_external_connection_export)       // external_connection.export
	);

	testbench_ls_input_IO input_io_1 (
		.clk        (clk_200_out_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_input_io_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_io_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_io_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_io_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_io_1_s1_readdata),   //                    .readdata
		.in_port    (input_io_1_external_connection_export)       // external_connection.export
	);

	testbench_ls_input_IO input_io_2 (
		.clk        (clk_200_out_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_input_io_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_io_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_io_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_io_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_io_2_s1_readdata),   //                    .readdata
		.in_port    (input_io_2_external_connection_export)       // external_connection.export
	);

	testbench_ls_input_IO input_io_3 (
		.clk        (clk_200_out_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_input_io_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_io_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_io_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_io_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_io_3_s1_readdata),   //                    .readdata
		.in_port    (input_io_3_external_connection_export)       // external_connection.export
	);

	testbench_ls_input_IO input_io_4 (
		.clk        (clk_200_out_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_input_io_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_io_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_io_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_io_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_io_4_s1_readdata),   //                    .readdata
		.in_port    (input_io_4_external_connection_export)       // external_connection.export
	);

	testbench_ls_input_IO_5 input_io_5 (
		.clk        (clk_200_out_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_input_io_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_io_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_io_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_io_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_io_5_s1_readdata),   //                    .readdata
		.in_port    (input_io_5_external_connection_export)       // external_connection.export
	);

	testbench_ls_jtag jtag (
		.clk            (clk_200_out_clk_clk),                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver6_irq)                              //               irq.irq
	);

	testbench_ls_nios_cpu nios_cpu (
		.clk                                 (clk_200_out_clk_clk),                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios_cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios_cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios_cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                        // custom_instruction_master.readra
	);

	testbench_ls_pilot_sig pilot_sig (
		.clk        (clk_200_out_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pilot_sig_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pilot_sig_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pilot_sig_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pilot_sig_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pilot_sig_s1_readdata),   //                    .readdata
		.in_port    (pilot_sig_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver8_irq)                   //                 irq.irq
	);

	testbench_ls_sys_timer sys_timer (
		.clk        (clk_200_out_clk_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_sys_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver7_irq)                   //   irq.irq
	);

	testbench_ls_system_ram system_ram (
		.clk        (clk_200_out_clk_clk),                        //   clk1.clk
		.address    (mm_interconnect_0_system_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_system_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_system_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_system_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_system_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_system_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_system_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	testbench_ls_mm_interconnect_0 mm_interconnect_0 (
		.ddr2_ram_afi_clk_clk                                        (clk_200_out_clk_clk),                                                     //                                      ddr2_ram_afi_clk.clk
		.ddr2_ram_1_afi_clk_clk                                      (ddr2_ram_1_afi_clk_clk),                                                  //                                    ddr2_ram_1_afi_clk.clk
		.ddr2_ram_1_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                                      // ddr2_ram_1_avl_translator_reset_reset_bridge_in_reset.reset
		.ddr2_ram_1_soft_reset_reset_bridge_in_reset_reset           (rst_controller_003_reset_out_reset),                                      //           ddr2_ram_1_soft_reset_reset_bridge_in_reset.reset
		.ddr2_ram_avl_translator_reset_reset_bridge_in_reset_reset   (rst_controller_004_reset_out_reset),                                      //   ddr2_ram_avl_translator_reset_reset_bridge_in_reset.reset
		.ddr2_ram_soft_reset_reset_bridge_in_reset_reset             (rst_controller_004_reset_out_reset),                                      //             ddr2_ram_soft_reset_reset_bridge_in_reset.reset
		.from_ETH_to_DDR_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                          //           from_ETH_to_DDR_reset_reset_bridge_in_reset.reset
		.nios_cpu_reset_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                                          //                  nios_cpu_reset_reset_bridge_in_reset.reset
		.dma_fifo_subsystem_1_dma_mm_read_address                    (dma_fifo_subsystem_1_dma_mm_read_address),                                //                      dma_fifo_subsystem_1_dma_mm_read.address
		.dma_fifo_subsystem_1_dma_mm_read_waitrequest                (dma_fifo_subsystem_1_dma_mm_read_waitrequest),                            //                                                      .waitrequest
		.dma_fifo_subsystem_1_dma_mm_read_burstcount                 (dma_fifo_subsystem_1_dma_mm_read_burstcount),                             //                                                      .burstcount
		.dma_fifo_subsystem_1_dma_mm_read_byteenable                 (dma_fifo_subsystem_1_dma_mm_read_byteenable),                             //                                                      .byteenable
		.dma_fifo_subsystem_1_dma_mm_read_read                       (dma_fifo_subsystem_1_dma_mm_read_read),                                   //                                                      .read
		.dma_fifo_subsystem_1_dma_mm_read_readdata                   (dma_fifo_subsystem_1_dma_mm_read_readdata),                               //                                                      .readdata
		.dma_fifo_subsystem_1_dma_mm_read_readdatavalid              (dma_fifo_subsystem_1_dma_mm_read_readdatavalid),                          //                                                      .readdatavalid
		.dma_fifo_subsystem_2_dma_mm_read_address                    (dma_fifo_subsystem_2_dma_mm_read_address),                                //                      dma_fifo_subsystem_2_dma_mm_read.address
		.dma_fifo_subsystem_2_dma_mm_read_waitrequest                (dma_fifo_subsystem_2_dma_mm_read_waitrequest),                            //                                                      .waitrequest
		.dma_fifo_subsystem_2_dma_mm_read_burstcount                 (dma_fifo_subsystem_2_dma_mm_read_burstcount),                             //                                                      .burstcount
		.dma_fifo_subsystem_2_dma_mm_read_byteenable                 (dma_fifo_subsystem_2_dma_mm_read_byteenable),                             //                                                      .byteenable
		.dma_fifo_subsystem_2_dma_mm_read_read                       (dma_fifo_subsystem_2_dma_mm_read_read),                                   //                                                      .read
		.dma_fifo_subsystem_2_dma_mm_read_readdata                   (dma_fifo_subsystem_2_dma_mm_read_readdata),                               //                                                      .readdata
		.dma_fifo_subsystem_2_dma_mm_read_readdatavalid              (dma_fifo_subsystem_2_dma_mm_read_readdatavalid),                          //                                                      .readdatavalid
		.dma_fifo_subsystem_3_dma_mm_read_address                    (dma_fifo_subsystem_3_dma_mm_read_address),                                //                      dma_fifo_subsystem_3_dma_mm_read.address
		.dma_fifo_subsystem_3_dma_mm_read_waitrequest                (dma_fifo_subsystem_3_dma_mm_read_waitrequest),                            //                                                      .waitrequest
		.dma_fifo_subsystem_3_dma_mm_read_burstcount                 (dma_fifo_subsystem_3_dma_mm_read_burstcount),                             //                                                      .burstcount
		.dma_fifo_subsystem_3_dma_mm_read_byteenable                 (dma_fifo_subsystem_3_dma_mm_read_byteenable),                             //                                                      .byteenable
		.dma_fifo_subsystem_3_dma_mm_read_read                       (dma_fifo_subsystem_3_dma_mm_read_read),                                   //                                                      .read
		.dma_fifo_subsystem_3_dma_mm_read_readdata                   (dma_fifo_subsystem_3_dma_mm_read_readdata),                               //                                                      .readdata
		.dma_fifo_subsystem_3_dma_mm_read_readdatavalid              (dma_fifo_subsystem_3_dma_mm_read_readdatavalid),                          //                                                      .readdatavalid
		.dma_fifo_subsystem_4_dma_mm_read_address                    (dma_fifo_subsystem_4_dma_mm_read_address),                                //                      dma_fifo_subsystem_4_dma_mm_read.address
		.dma_fifo_subsystem_4_dma_mm_read_waitrequest                (dma_fifo_subsystem_4_dma_mm_read_waitrequest),                            //                                                      .waitrequest
		.dma_fifo_subsystem_4_dma_mm_read_burstcount                 (dma_fifo_subsystem_4_dma_mm_read_burstcount),                             //                                                      .burstcount
		.dma_fifo_subsystem_4_dma_mm_read_byteenable                 (dma_fifo_subsystem_4_dma_mm_read_byteenable),                             //                                                      .byteenable
		.dma_fifo_subsystem_4_dma_mm_read_read                       (dma_fifo_subsystem_4_dma_mm_read_read),                                   //                                                      .read
		.dma_fifo_subsystem_4_dma_mm_read_readdata                   (dma_fifo_subsystem_4_dma_mm_read_readdata),                               //                                                      .readdata
		.dma_fifo_subsystem_4_dma_mm_read_readdatavalid              (dma_fifo_subsystem_4_dma_mm_read_readdatavalid),                          //                                                      .readdatavalid
		.dma_fifo_susbystem_dma_mm_read_address                      (dma_fifo_susbystem_dma_mm_read_address),                                  //                        dma_fifo_susbystem_dma_mm_read.address
		.dma_fifo_susbystem_dma_mm_read_waitrequest                  (dma_fifo_susbystem_dma_mm_read_waitrequest),                              //                                                      .waitrequest
		.dma_fifo_susbystem_dma_mm_read_burstcount                   (dma_fifo_susbystem_dma_mm_read_burstcount),                               //                                                      .burstcount
		.dma_fifo_susbystem_dma_mm_read_byteenable                   (dma_fifo_susbystem_dma_mm_read_byteenable),                               //                                                      .byteenable
		.dma_fifo_susbystem_dma_mm_read_read                         (dma_fifo_susbystem_dma_mm_read_read),                                     //                                                      .read
		.dma_fifo_susbystem_dma_mm_read_readdata                     (dma_fifo_susbystem_dma_mm_read_readdata),                                 //                                                      .readdata
		.dma_fifo_susbystem_dma_mm_read_readdatavalid                (dma_fifo_susbystem_dma_mm_read_readdatavalid),                            //                                                      .readdatavalid
		.from_ETH_to_DDR_ETH_DMA_mm_write_address                    (from_eth_to_ddr_eth_dma_mm_write_address),                                //                      from_ETH_to_DDR_ETH_DMA_mm_write.address
		.from_ETH_to_DDR_ETH_DMA_mm_write_waitrequest                (from_eth_to_ddr_eth_dma_mm_write_waitrequest),                            //                                                      .waitrequest
		.from_ETH_to_DDR_ETH_DMA_mm_write_byteenable                 (from_eth_to_ddr_eth_dma_mm_write_byteenable),                             //                                                      .byteenable
		.from_ETH_to_DDR_ETH_DMA_mm_write_write                      (from_eth_to_ddr_eth_dma_mm_write_write),                                  //                                                      .write
		.from_ETH_to_DDR_ETH_DMA_mm_write_writedata                  (from_eth_to_ddr_eth_dma_mm_write_writedata),                              //                                                      .writedata
		.nios_cpu_data_master_address                                (nios_cpu_data_master_address),                                            //                                  nios_cpu_data_master.address
		.nios_cpu_data_master_waitrequest                            (nios_cpu_data_master_waitrequest),                                        //                                                      .waitrequest
		.nios_cpu_data_master_byteenable                             (nios_cpu_data_master_byteenable),                                         //                                                      .byteenable
		.nios_cpu_data_master_read                                   (nios_cpu_data_master_read),                                               //                                                      .read
		.nios_cpu_data_master_readdata                               (nios_cpu_data_master_readdata),                                           //                                                      .readdata
		.nios_cpu_data_master_readdatavalid                          (nios_cpu_data_master_readdatavalid),                                      //                                                      .readdatavalid
		.nios_cpu_data_master_write                                  (nios_cpu_data_master_write),                                              //                                                      .write
		.nios_cpu_data_master_writedata                              (nios_cpu_data_master_writedata),                                          //                                                      .writedata
		.nios_cpu_data_master_debugaccess                            (nios_cpu_data_master_debugaccess),                                        //                                                      .debugaccess
		.nios_cpu_instruction_master_address                         (nios_cpu_instruction_master_address),                                     //                           nios_cpu_instruction_master.address
		.nios_cpu_instruction_master_waitrequest                     (nios_cpu_instruction_master_waitrequest),                                 //                                                      .waitrequest
		.nios_cpu_instruction_master_read                            (nios_cpu_instruction_master_read),                                        //                                                      .read
		.nios_cpu_instruction_master_readdata                        (nios_cpu_instruction_master_readdata),                                    //                                                      .readdata
		.nios_cpu_instruction_master_readdatavalid                   (nios_cpu_instruction_master_readdatavalid),                               //                                                      .readdatavalid
		.ctrl_sig_s1_address                                         (mm_interconnect_0_ctrl_sig_s1_address),                                   //                                           ctrl_sig_s1.address
		.ctrl_sig_s1_write                                           (mm_interconnect_0_ctrl_sig_s1_write),                                     //                                                      .write
		.ctrl_sig_s1_readdata                                        (mm_interconnect_0_ctrl_sig_s1_readdata),                                  //                                                      .readdata
		.ctrl_sig_s1_writedata                                       (mm_interconnect_0_ctrl_sig_s1_writedata),                                 //                                                      .writedata
		.ctrl_sig_s1_chipselect                                      (mm_interconnect_0_ctrl_sig_s1_chipselect),                                //                                                      .chipselect
		.ddr2_ram_avl_address                                        (mm_interconnect_0_ddr2_ram_avl_address),                                  //                                          ddr2_ram_avl.address
		.ddr2_ram_avl_write                                          (mm_interconnect_0_ddr2_ram_avl_write),                                    //                                                      .write
		.ddr2_ram_avl_read                                           (mm_interconnect_0_ddr2_ram_avl_read),                                     //                                                      .read
		.ddr2_ram_avl_readdata                                       (mm_interconnect_0_ddr2_ram_avl_readdata),                                 //                                                      .readdata
		.ddr2_ram_avl_writedata                                      (mm_interconnect_0_ddr2_ram_avl_writedata),                                //                                                      .writedata
		.ddr2_ram_avl_beginbursttransfer                             (mm_interconnect_0_ddr2_ram_avl_beginbursttransfer),                       //                                                      .beginbursttransfer
		.ddr2_ram_avl_burstcount                                     (mm_interconnect_0_ddr2_ram_avl_burstcount),                               //                                                      .burstcount
		.ddr2_ram_avl_byteenable                                     (mm_interconnect_0_ddr2_ram_avl_byteenable),                               //                                                      .byteenable
		.ddr2_ram_avl_readdatavalid                                  (mm_interconnect_0_ddr2_ram_avl_readdatavalid),                            //                                                      .readdatavalid
		.ddr2_ram_avl_waitrequest                                    (~mm_interconnect_0_ddr2_ram_avl_waitrequest),                             //                                                      .waitrequest
		.ddr2_ram_1_avl_address                                      (mm_interconnect_0_ddr2_ram_1_avl_address),                                //                                        ddr2_ram_1_avl.address
		.ddr2_ram_1_avl_write                                        (mm_interconnect_0_ddr2_ram_1_avl_write),                                  //                                                      .write
		.ddr2_ram_1_avl_read                                         (mm_interconnect_0_ddr2_ram_1_avl_read),                                   //                                                      .read
		.ddr2_ram_1_avl_readdata                                     (mm_interconnect_0_ddr2_ram_1_avl_readdata),                               //                                                      .readdata
		.ddr2_ram_1_avl_writedata                                    (mm_interconnect_0_ddr2_ram_1_avl_writedata),                              //                                                      .writedata
		.ddr2_ram_1_avl_beginbursttransfer                           (mm_interconnect_0_ddr2_ram_1_avl_beginbursttransfer),                     //                                                      .beginbursttransfer
		.ddr2_ram_1_avl_burstcount                                   (mm_interconnect_0_ddr2_ram_1_avl_burstcount),                             //                                                      .burstcount
		.ddr2_ram_1_avl_byteenable                                   (mm_interconnect_0_ddr2_ram_1_avl_byteenable),                             //                                                      .byteenable
		.ddr2_ram_1_avl_readdatavalid                                (mm_interconnect_0_ddr2_ram_1_avl_readdatavalid),                          //                                                      .readdatavalid
		.ddr2_ram_1_avl_waitrequest                                  (~mm_interconnect_0_ddr2_ram_1_avl_waitrequest),                           //                                                      .waitrequest
		.dma_fifo_subsystem_1_dma_csr_address                        (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_address),                  //                          dma_fifo_subsystem_1_dma_csr.address
		.dma_fifo_subsystem_1_dma_csr_write                          (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_write),                    //                                                      .write
		.dma_fifo_subsystem_1_dma_csr_read                           (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_read),                     //                                                      .read
		.dma_fifo_subsystem_1_dma_csr_readdata                       (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_readdata),                 //                                                      .readdata
		.dma_fifo_subsystem_1_dma_csr_writedata                      (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_writedata),                //                                                      .writedata
		.dma_fifo_subsystem_1_dma_csr_byteenable                     (mm_interconnect_0_dma_fifo_subsystem_1_dma_csr_byteenable),               //                                                      .byteenable
		.dma_fifo_subsystem_1_dma_descriptor_slave_write             (mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_write),       //             dma_fifo_subsystem_1_dma_descriptor_slave.write
		.dma_fifo_subsystem_1_dma_descriptor_slave_writedata         (mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_writedata),   //                                                      .writedata
		.dma_fifo_subsystem_1_dma_descriptor_slave_byteenable        (mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_byteenable),  //                                                      .byteenable
		.dma_fifo_subsystem_1_dma_descriptor_slave_waitrequest       (mm_interconnect_0_dma_fifo_subsystem_1_dma_descriptor_slave_waitrequest), //                                                      .waitrequest
		.dma_fifo_subsystem_2_dma_csr_address                        (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_address),                  //                          dma_fifo_subsystem_2_dma_csr.address
		.dma_fifo_subsystem_2_dma_csr_write                          (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_write),                    //                                                      .write
		.dma_fifo_subsystem_2_dma_csr_read                           (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_read),                     //                                                      .read
		.dma_fifo_subsystem_2_dma_csr_readdata                       (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_readdata),                 //                                                      .readdata
		.dma_fifo_subsystem_2_dma_csr_writedata                      (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_writedata),                //                                                      .writedata
		.dma_fifo_subsystem_2_dma_csr_byteenable                     (mm_interconnect_0_dma_fifo_subsystem_2_dma_csr_byteenable),               //                                                      .byteenable
		.dma_fifo_subsystem_2_dma_descriptor_slave_write             (mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_write),       //             dma_fifo_subsystem_2_dma_descriptor_slave.write
		.dma_fifo_subsystem_2_dma_descriptor_slave_writedata         (mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_writedata),   //                                                      .writedata
		.dma_fifo_subsystem_2_dma_descriptor_slave_byteenable        (mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_byteenable),  //                                                      .byteenable
		.dma_fifo_subsystem_2_dma_descriptor_slave_waitrequest       (mm_interconnect_0_dma_fifo_subsystem_2_dma_descriptor_slave_waitrequest), //                                                      .waitrequest
		.dma_fifo_subsystem_3_dma_csr_address                        (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_address),                  //                          dma_fifo_subsystem_3_dma_csr.address
		.dma_fifo_subsystem_3_dma_csr_write                          (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_write),                    //                                                      .write
		.dma_fifo_subsystem_3_dma_csr_read                           (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_read),                     //                                                      .read
		.dma_fifo_subsystem_3_dma_csr_readdata                       (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_readdata),                 //                                                      .readdata
		.dma_fifo_subsystem_3_dma_csr_writedata                      (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_writedata),                //                                                      .writedata
		.dma_fifo_subsystem_3_dma_csr_byteenable                     (mm_interconnect_0_dma_fifo_subsystem_3_dma_csr_byteenable),               //                                                      .byteenable
		.dma_fifo_subsystem_3_dma_descriptor_slave_write             (mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_write),       //             dma_fifo_subsystem_3_dma_descriptor_slave.write
		.dma_fifo_subsystem_3_dma_descriptor_slave_writedata         (mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_writedata),   //                                                      .writedata
		.dma_fifo_subsystem_3_dma_descriptor_slave_byteenable        (mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_byteenable),  //                                                      .byteenable
		.dma_fifo_subsystem_3_dma_descriptor_slave_waitrequest       (mm_interconnect_0_dma_fifo_subsystem_3_dma_descriptor_slave_waitrequest), //                                                      .waitrequest
		.dma_fifo_subsystem_4_dma_csr_address                        (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_address),                  //                          dma_fifo_subsystem_4_dma_csr.address
		.dma_fifo_subsystem_4_dma_csr_write                          (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_write),                    //                                                      .write
		.dma_fifo_subsystem_4_dma_csr_read                           (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_read),                     //                                                      .read
		.dma_fifo_subsystem_4_dma_csr_readdata                       (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_readdata),                 //                                                      .readdata
		.dma_fifo_subsystem_4_dma_csr_writedata                      (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_writedata),                //                                                      .writedata
		.dma_fifo_subsystem_4_dma_csr_byteenable                     (mm_interconnect_0_dma_fifo_subsystem_4_dma_csr_byteenable),               //                                                      .byteenable
		.dma_fifo_subsystem_4_dma_descriptor_slave_write             (mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_write),       //             dma_fifo_subsystem_4_dma_descriptor_slave.write
		.dma_fifo_subsystem_4_dma_descriptor_slave_writedata         (mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_writedata),   //                                                      .writedata
		.dma_fifo_subsystem_4_dma_descriptor_slave_byteenable        (mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_byteenable),  //                                                      .byteenable
		.dma_fifo_subsystem_4_dma_descriptor_slave_waitrequest       (mm_interconnect_0_dma_fifo_subsystem_4_dma_descriptor_slave_waitrequest), //                                                      .waitrequest
		.dma_fifo_susbystem_dma_csr_address                          (mm_interconnect_0_dma_fifo_susbystem_dma_csr_address),                    //                            dma_fifo_susbystem_dma_csr.address
		.dma_fifo_susbystem_dma_csr_write                            (mm_interconnect_0_dma_fifo_susbystem_dma_csr_write),                      //                                                      .write
		.dma_fifo_susbystem_dma_csr_read                             (mm_interconnect_0_dma_fifo_susbystem_dma_csr_read),                       //                                                      .read
		.dma_fifo_susbystem_dma_csr_readdata                         (mm_interconnect_0_dma_fifo_susbystem_dma_csr_readdata),                   //                                                      .readdata
		.dma_fifo_susbystem_dma_csr_writedata                        (mm_interconnect_0_dma_fifo_susbystem_dma_csr_writedata),                  //                                                      .writedata
		.dma_fifo_susbystem_dma_csr_byteenable                       (mm_interconnect_0_dma_fifo_susbystem_dma_csr_byteenable),                 //                                                      .byteenable
		.dma_fifo_susbystem_dma_descriptor_slave_write               (mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_write),         //               dma_fifo_susbystem_dma_descriptor_slave.write
		.dma_fifo_susbystem_dma_descriptor_slave_writedata           (mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_writedata),     //                                                      .writedata
		.dma_fifo_susbystem_dma_descriptor_slave_byteenable          (mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_byteenable),    //                                                      .byteenable
		.dma_fifo_susbystem_dma_descriptor_slave_waitrequest         (mm_interconnect_0_dma_fifo_susbystem_dma_descriptor_slave_waitrequest),   //                                                      .waitrequest
		.from_ETH_to_DDR_ETH_DMA_csr_address                         (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_address),                   //                           from_ETH_to_DDR_ETH_DMA_csr.address
		.from_ETH_to_DDR_ETH_DMA_csr_write                           (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_write),                     //                                                      .write
		.from_ETH_to_DDR_ETH_DMA_csr_read                            (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_read),                      //                                                      .read
		.from_ETH_to_DDR_ETH_DMA_csr_readdata                        (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_readdata),                  //                                                      .readdata
		.from_ETH_to_DDR_ETH_DMA_csr_writedata                       (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_writedata),                 //                                                      .writedata
		.from_ETH_to_DDR_ETH_DMA_csr_byteenable                      (mm_interconnect_0_from_eth_to_ddr_eth_dma_csr_byteenable),                //                                                      .byteenable
		.from_ETH_to_DDR_ETH_DMA_descriptor_slave_write              (mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_write),        //              from_ETH_to_DDR_ETH_DMA_descriptor_slave.write
		.from_ETH_to_DDR_ETH_DMA_descriptor_slave_writedata          (mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_writedata),    //                                                      .writedata
		.from_ETH_to_DDR_ETH_DMA_descriptor_slave_byteenable         (mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_byteenable),   //                                                      .byteenable
		.from_ETH_to_DDR_ETH_DMA_descriptor_slave_waitrequest        (mm_interconnect_0_from_eth_to_ddr_eth_dma_descriptor_slave_waitrequest),  //                                                      .waitrequest
		.input_IO_s1_address                                         (mm_interconnect_0_input_io_s1_address),                                   //                                           input_IO_s1.address
		.input_IO_s1_write                                           (mm_interconnect_0_input_io_s1_write),                                     //                                                      .write
		.input_IO_s1_readdata                                        (mm_interconnect_0_input_io_s1_readdata),                                  //                                                      .readdata
		.input_IO_s1_writedata                                       (mm_interconnect_0_input_io_s1_writedata),                                 //                                                      .writedata
		.input_IO_s1_chipselect                                      (mm_interconnect_0_input_io_s1_chipselect),                                //                                                      .chipselect
		.input_IO_0_s1_address                                       (mm_interconnect_0_input_io_0_s1_address),                                 //                                         input_IO_0_s1.address
		.input_IO_0_s1_write                                         (mm_interconnect_0_input_io_0_s1_write),                                   //                                                      .write
		.input_IO_0_s1_readdata                                      (mm_interconnect_0_input_io_0_s1_readdata),                                //                                                      .readdata
		.input_IO_0_s1_writedata                                     (mm_interconnect_0_input_io_0_s1_writedata),                               //                                                      .writedata
		.input_IO_0_s1_chipselect                                    (mm_interconnect_0_input_io_0_s1_chipselect),                              //                                                      .chipselect
		.input_IO_1_s1_address                                       (mm_interconnect_0_input_io_1_s1_address),                                 //                                         input_IO_1_s1.address
		.input_IO_1_s1_write                                         (mm_interconnect_0_input_io_1_s1_write),                                   //                                                      .write
		.input_IO_1_s1_readdata                                      (mm_interconnect_0_input_io_1_s1_readdata),                                //                                                      .readdata
		.input_IO_1_s1_writedata                                     (mm_interconnect_0_input_io_1_s1_writedata),                               //                                                      .writedata
		.input_IO_1_s1_chipselect                                    (mm_interconnect_0_input_io_1_s1_chipselect),                              //                                                      .chipselect
		.input_IO_2_s1_address                                       (mm_interconnect_0_input_io_2_s1_address),                                 //                                         input_IO_2_s1.address
		.input_IO_2_s1_write                                         (mm_interconnect_0_input_io_2_s1_write),                                   //                                                      .write
		.input_IO_2_s1_readdata                                      (mm_interconnect_0_input_io_2_s1_readdata),                                //                                                      .readdata
		.input_IO_2_s1_writedata                                     (mm_interconnect_0_input_io_2_s1_writedata),                               //                                                      .writedata
		.input_IO_2_s1_chipselect                                    (mm_interconnect_0_input_io_2_s1_chipselect),                              //                                                      .chipselect
		.input_IO_3_s1_address                                       (mm_interconnect_0_input_io_3_s1_address),                                 //                                         input_IO_3_s1.address
		.input_IO_3_s1_write                                         (mm_interconnect_0_input_io_3_s1_write),                                   //                                                      .write
		.input_IO_3_s1_readdata                                      (mm_interconnect_0_input_io_3_s1_readdata),                                //                                                      .readdata
		.input_IO_3_s1_writedata                                     (mm_interconnect_0_input_io_3_s1_writedata),                               //                                                      .writedata
		.input_IO_3_s1_chipselect                                    (mm_interconnect_0_input_io_3_s1_chipselect),                              //                                                      .chipselect
		.input_IO_4_s1_address                                       (mm_interconnect_0_input_io_4_s1_address),                                 //                                         input_IO_4_s1.address
		.input_IO_4_s1_write                                         (mm_interconnect_0_input_io_4_s1_write),                                   //                                                      .write
		.input_IO_4_s1_readdata                                      (mm_interconnect_0_input_io_4_s1_readdata),                                //                                                      .readdata
		.input_IO_4_s1_writedata                                     (mm_interconnect_0_input_io_4_s1_writedata),                               //                                                      .writedata
		.input_IO_4_s1_chipselect                                    (mm_interconnect_0_input_io_4_s1_chipselect),                              //                                                      .chipselect
		.input_IO_5_s1_address                                       (mm_interconnect_0_input_io_5_s1_address),                                 //                                         input_IO_5_s1.address
		.input_IO_5_s1_write                                         (mm_interconnect_0_input_io_5_s1_write),                                   //                                                      .write
		.input_IO_5_s1_readdata                                      (mm_interconnect_0_input_io_5_s1_readdata),                                //                                                      .readdata
		.input_IO_5_s1_writedata                                     (mm_interconnect_0_input_io_5_s1_writedata),                               //                                                      .writedata
		.input_IO_5_s1_chipselect                                    (mm_interconnect_0_input_io_5_s1_chipselect),                              //                                                      .chipselect
		.jtag_avalon_jtag_slave_address                              (mm_interconnect_0_jtag_avalon_jtag_slave_address),                        //                                jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                                (mm_interconnect_0_jtag_avalon_jtag_slave_write),                          //                                                      .write
		.jtag_avalon_jtag_slave_read                                 (mm_interconnect_0_jtag_avalon_jtag_slave_read),                           //                                                      .read
		.jtag_avalon_jtag_slave_readdata                             (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                       //                                                      .readdata
		.jtag_avalon_jtag_slave_writedata                            (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),                      //                                                      .writedata
		.jtag_avalon_jtag_slave_waitrequest                          (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),                    //                                                      .waitrequest
		.jtag_avalon_jtag_slave_chipselect                           (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),                     //                                                      .chipselect
		.nios_cpu_debug_mem_slave_address                            (mm_interconnect_0_nios_cpu_debug_mem_slave_address),                      //                              nios_cpu_debug_mem_slave.address
		.nios_cpu_debug_mem_slave_write                              (mm_interconnect_0_nios_cpu_debug_mem_slave_write),                        //                                                      .write
		.nios_cpu_debug_mem_slave_read                               (mm_interconnect_0_nios_cpu_debug_mem_slave_read),                         //                                                      .read
		.nios_cpu_debug_mem_slave_readdata                           (mm_interconnect_0_nios_cpu_debug_mem_slave_readdata),                     //                                                      .readdata
		.nios_cpu_debug_mem_slave_writedata                          (mm_interconnect_0_nios_cpu_debug_mem_slave_writedata),                    //                                                      .writedata
		.nios_cpu_debug_mem_slave_byteenable                         (mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable),                   //                                                      .byteenable
		.nios_cpu_debug_mem_slave_waitrequest                        (mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest),                  //                                                      .waitrequest
		.nios_cpu_debug_mem_slave_debugaccess                        (mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess),                  //                                                      .debugaccess
		.pilot_sig_s1_address                                        (mm_interconnect_0_pilot_sig_s1_address),                                  //                                          pilot_sig_s1.address
		.pilot_sig_s1_write                                          (mm_interconnect_0_pilot_sig_s1_write),                                    //                                                      .write
		.pilot_sig_s1_readdata                                       (mm_interconnect_0_pilot_sig_s1_readdata),                                 //                                                      .readdata
		.pilot_sig_s1_writedata                                      (mm_interconnect_0_pilot_sig_s1_writedata),                                //                                                      .writedata
		.pilot_sig_s1_chipselect                                     (mm_interconnect_0_pilot_sig_s1_chipselect),                               //                                                      .chipselect
		.sys_timer_s1_address                                        (mm_interconnect_0_sys_timer_s1_address),                                  //                                          sys_timer_s1.address
		.sys_timer_s1_write                                          (mm_interconnect_0_sys_timer_s1_write),                                    //                                                      .write
		.sys_timer_s1_readdata                                       (mm_interconnect_0_sys_timer_s1_readdata),                                 //                                                      .readdata
		.sys_timer_s1_writedata                                      (mm_interconnect_0_sys_timer_s1_writedata),                                //                                                      .writedata
		.sys_timer_s1_chipselect                                     (mm_interconnect_0_sys_timer_s1_chipselect),                               //                                                      .chipselect
		.system_ram_s1_address                                       (mm_interconnect_0_system_ram_s1_address),                                 //                                         system_ram_s1.address
		.system_ram_s1_write                                         (mm_interconnect_0_system_ram_s1_write),                                   //                                                      .write
		.system_ram_s1_readdata                                      (mm_interconnect_0_system_ram_s1_readdata),                                //                                                      .readdata
		.system_ram_s1_writedata                                     (mm_interconnect_0_system_ram_s1_writedata),                               //                                                      .writedata
		.system_ram_s1_byteenable                                    (mm_interconnect_0_system_ram_s1_byteenable),                              //                                                      .byteenable
		.system_ram_s1_chipselect                                    (mm_interconnect_0_system_ram_s1_chipselect),                              //                                                      .chipselect
		.system_ram_s1_clken                                         (mm_interconnect_0_system_ram_s1_clken)                                    //                                                      .clken
	);

	testbench_ls_irq_mapper irq_mapper (
		.clk           (clk_200_out_clk_clk),            //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),       // receiver8.irq
		.sender_irq    (nios_cpu_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_200_out_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (ddr2_ram_1_afi_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_200_out_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
